VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_w6_r100
  CLASS BLOCK ;
  FOREIGN vco_w6_r100 ;
  ORIGIN 0.450 12.000 ;
  SIZE 123.580 BY 105.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 92.420 33.250 92.800 33.300 ;
        RECT 91.470 32.890 92.800 33.250 ;
        RECT 92.420 32.840 92.800 32.890 ;
        RECT 94.290 33.250 94.670 33.300 ;
        RECT 94.290 32.890 95.620 33.250 ;
        RECT 94.290 32.840 94.670 32.890 ;
        RECT 96.730 26.750 97.030 39.340 ;
        RECT 100.960 33.250 101.340 33.300 ;
        RECT 100.960 32.890 102.290 33.250 ;
        RECT 100.960 32.840 101.340 32.890 ;
        RECT 111.105 26.750 111.405 39.340 ;
      LAYER mcon ;
        RECT 91.470 32.920 91.770 33.220 ;
        RECT 91.960 32.920 92.260 33.220 ;
        RECT 92.450 32.920 92.750 33.220 ;
        RECT 94.340 32.920 94.640 33.220 ;
        RECT 94.830 32.920 95.130 33.220 ;
        RECT 95.320 32.920 95.620 33.220 ;
        RECT 101.010 32.920 101.310 33.220 ;
        RECT 101.500 32.920 101.800 33.220 ;
        RECT 101.990 32.920 102.290 33.220 ;
        RECT 96.730 31.560 97.030 31.860 ;
        RECT 111.105 31.560 111.405 31.860 ;
      LAYER met1 ;
        RECT 91.410 32.890 95.680 33.250 ;
        RECT 100.850 32.890 102.350 33.250 ;
        RECT 94.710 31.890 95.070 32.890 ;
        RECT 101.440 31.890 101.800 32.890 ;
        RECT 94.710 31.530 111.465 31.890 ;
      LAYER via ;
        RECT 96.140 31.530 96.500 31.890 ;
      LAYER met2 ;
        RECT 96.110 24.280 96.530 31.890 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 74.710 33.250 75.090 33.300 ;
        RECT 73.760 32.890 75.090 33.250 ;
        RECT 74.710 32.840 75.090 32.890 ;
        RECT 76.580 33.250 76.960 33.300 ;
        RECT 76.580 32.890 77.910 33.250 ;
        RECT 76.580 32.840 76.960 32.890 ;
        RECT 79.020 26.750 79.320 39.340 ;
        RECT 83.250 33.250 83.630 33.300 ;
        RECT 83.250 32.890 84.580 33.250 ;
        RECT 83.250 32.840 83.630 32.890 ;
        RECT 93.395 26.750 93.695 39.340 ;
      LAYER mcon ;
        RECT 73.760 32.920 74.060 33.220 ;
        RECT 74.250 32.920 74.550 33.220 ;
        RECT 74.740 32.920 75.040 33.220 ;
        RECT 76.630 32.920 76.930 33.220 ;
        RECT 77.120 32.920 77.420 33.220 ;
        RECT 77.610 32.920 77.910 33.220 ;
        RECT 83.300 32.920 83.600 33.220 ;
        RECT 83.790 32.920 84.090 33.220 ;
        RECT 84.280 32.920 84.580 33.220 ;
        RECT 79.020 31.560 79.320 31.860 ;
        RECT 93.395 31.560 93.695 31.860 ;
      LAYER met1 ;
        RECT 73.700 32.890 77.970 33.250 ;
        RECT 83.140 32.890 84.640 33.250 ;
        RECT 77.000 31.890 77.360 32.890 ;
        RECT 83.730 31.890 84.090 32.890 ;
        RECT 77.000 31.530 93.755 31.890 ;
      LAYER via ;
        RECT 79.340 31.530 79.700 31.890 ;
      LAYER met2 ;
        RECT 79.310 24.280 79.730 31.890 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 57.000 33.250 57.380 33.300 ;
        RECT 56.050 32.890 57.380 33.250 ;
        RECT 57.000 32.840 57.380 32.890 ;
        RECT 58.870 33.250 59.250 33.300 ;
        RECT 58.870 32.890 60.200 33.250 ;
        RECT 58.870 32.840 59.250 32.890 ;
        RECT 61.310 26.750 61.610 39.340 ;
        RECT 65.540 33.250 65.920 33.300 ;
        RECT 65.540 32.890 66.870 33.250 ;
        RECT 65.540 32.840 65.920 32.890 ;
        RECT 75.685 26.750 75.985 39.340 ;
      LAYER mcon ;
        RECT 56.050 32.920 56.350 33.220 ;
        RECT 56.540 32.920 56.840 33.220 ;
        RECT 57.030 32.920 57.330 33.220 ;
        RECT 58.920 32.920 59.220 33.220 ;
        RECT 59.410 32.920 59.710 33.220 ;
        RECT 59.900 32.920 60.200 33.220 ;
        RECT 65.590 32.920 65.890 33.220 ;
        RECT 66.080 32.920 66.380 33.220 ;
        RECT 66.570 32.920 66.870 33.220 ;
        RECT 61.310 31.560 61.610 31.860 ;
        RECT 75.685 31.560 75.985 31.860 ;
      LAYER met1 ;
        RECT 55.990 32.890 60.260 33.250 ;
        RECT 65.430 32.890 66.930 33.250 ;
        RECT 59.290 31.890 59.650 32.890 ;
        RECT 66.020 31.890 66.380 32.890 ;
        RECT 59.290 31.530 76.045 31.890 ;
      LAYER via ;
        RECT 66.020 31.530 66.380 31.890 ;
      LAYER met2 ;
        RECT 65.990 24.280 66.410 31.890 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 39.290 33.250 39.670 33.300 ;
        RECT 38.340 32.890 39.670 33.250 ;
        RECT 39.290 32.840 39.670 32.890 ;
        RECT 41.160 33.250 41.540 33.300 ;
        RECT 41.160 32.890 42.490 33.250 ;
        RECT 41.160 32.840 41.540 32.890 ;
        RECT 43.600 26.750 43.900 39.340 ;
        RECT 47.830 33.250 48.210 33.300 ;
        RECT 47.830 32.890 49.160 33.250 ;
        RECT 47.830 32.840 48.210 32.890 ;
        RECT 57.975 26.750 58.275 39.340 ;
      LAYER mcon ;
        RECT 38.340 32.920 38.640 33.220 ;
        RECT 38.830 32.920 39.130 33.220 ;
        RECT 39.320 32.920 39.620 33.220 ;
        RECT 41.210 32.920 41.510 33.220 ;
        RECT 41.700 32.920 42.000 33.220 ;
        RECT 42.190 32.920 42.490 33.220 ;
        RECT 47.880 32.920 48.180 33.220 ;
        RECT 48.370 32.920 48.670 33.220 ;
        RECT 48.860 32.920 49.160 33.220 ;
        RECT 43.600 31.560 43.900 31.860 ;
        RECT 57.975 31.560 58.275 31.860 ;
      LAYER met1 ;
        RECT 38.280 32.890 42.550 33.250 ;
        RECT 47.720 32.890 49.220 33.250 ;
        RECT 41.580 31.890 41.940 32.890 ;
        RECT 48.310 31.890 48.670 32.890 ;
        RECT 41.580 31.530 58.335 31.890 ;
      LAYER via ;
        RECT 43.030 31.530 43.390 31.890 ;
      LAYER met2 ;
        RECT 43.000 24.280 43.420 31.890 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 21.580 33.250 21.960 33.300 ;
        RECT 20.630 32.890 21.960 33.250 ;
        RECT 21.580 32.840 21.960 32.890 ;
        RECT 23.450 33.250 23.830 33.300 ;
        RECT 23.450 32.890 24.780 33.250 ;
        RECT 23.450 32.840 23.830 32.890 ;
        RECT 25.890 26.750 26.190 39.340 ;
        RECT 30.120 33.250 30.500 33.300 ;
        RECT 30.120 32.890 31.450 33.250 ;
        RECT 30.120 32.840 30.500 32.890 ;
        RECT 40.265 26.750 40.565 39.340 ;
      LAYER mcon ;
        RECT 20.630 32.920 20.930 33.220 ;
        RECT 21.120 32.920 21.420 33.220 ;
        RECT 21.610 32.920 21.910 33.220 ;
        RECT 23.500 32.920 23.800 33.220 ;
        RECT 23.990 32.920 24.290 33.220 ;
        RECT 24.480 32.920 24.780 33.220 ;
        RECT 30.170 32.920 30.470 33.220 ;
        RECT 30.660 32.920 30.960 33.220 ;
        RECT 31.150 32.920 31.450 33.220 ;
        RECT 25.890 31.560 26.190 31.860 ;
        RECT 40.265 31.560 40.565 31.860 ;
      LAYER met1 ;
        RECT 20.570 32.890 24.840 33.250 ;
        RECT 30.010 32.890 31.510 33.250 ;
        RECT 23.870 31.890 24.230 32.890 ;
        RECT 30.600 31.890 30.960 32.890 ;
        RECT 23.870 31.530 40.625 31.890 ;
      LAYER via ;
        RECT 25.280 31.530 25.640 31.890 ;
      LAYER met2 ;
        RECT 25.250 24.280 25.670 31.890 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 6.245500 ;
    PORT
      LAYER li1 ;
        RECT 8.310 50.925 8.905 51.265 ;
        RECT 8.310 49.605 8.485 50.925 ;
        RECT 8.310 49.480 8.905 49.605 ;
        RECT 9.710 49.480 10.010 50.310 ;
        RECT 8.310 49.180 10.010 49.480 ;
        RECT 8.310 49.055 8.905 49.180 ;
        RECT 17.880 48.950 18.260 49.000 ;
        RECT 16.930 48.590 18.260 48.950 ;
        RECT 17.880 48.540 18.260 48.590 ;
        RECT 19.750 48.950 20.130 49.000 ;
        RECT 19.750 48.590 21.080 48.950 ;
        RECT 19.750 48.540 20.130 48.590 ;
        RECT 8.180 26.750 8.480 39.340 ;
        RECT 12.410 33.250 12.790 33.300 ;
        RECT 12.410 32.890 13.740 33.250 ;
        RECT 12.410 32.840 12.790 32.890 ;
        RECT 22.555 26.750 22.855 39.340 ;
      LAYER mcon ;
        RECT 9.740 50.040 9.980 50.280 ;
        RECT 16.930 48.620 17.230 48.920 ;
        RECT 17.420 48.620 17.720 48.920 ;
        RECT 17.910 48.620 18.210 48.920 ;
        RECT 19.800 48.620 20.100 48.920 ;
        RECT 20.290 48.620 20.590 48.920 ;
        RECT 20.780 48.620 21.080 48.920 ;
        RECT 12.460 32.920 12.760 33.220 ;
        RECT 12.950 32.920 13.250 33.220 ;
        RECT 13.440 32.920 13.740 33.220 ;
        RECT 8.180 31.560 8.480 31.860 ;
        RECT 22.555 31.560 22.855 31.860 ;
      LAYER met1 ;
        RECT 9.680 50.010 17.840 50.310 ;
        RECT 13.260 49.950 17.840 50.010 ;
        RECT 13.260 43.360 13.620 49.950 ;
        RECT 17.480 48.950 17.840 49.950 ;
        RECT 16.870 48.590 21.140 48.950 ;
        RECT 4.990 43.000 13.620 43.360 ;
        RECT 4.990 31.890 5.350 43.000 ;
        RECT 12.300 32.890 13.800 33.250 ;
        RECT 12.890 31.890 13.250 32.890 ;
        RECT 4.990 31.530 22.915 31.890 ;
      LAYER via ;
        RECT 7.140 31.530 7.500 31.890 ;
      LAYER met2 ;
        RECT 7.110 24.280 7.530 31.890 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 18.855 42.500 19.155 55.090 ;
        RECT 28.920 48.950 29.300 49.000 ;
        RECT 27.970 48.590 29.300 48.950 ;
        RECT 28.920 48.540 29.300 48.590 ;
        RECT 33.230 42.500 33.530 55.090 ;
        RECT 35.590 48.950 35.970 49.000 ;
        RECT 34.640 48.590 35.970 48.950 ;
        RECT 35.590 48.540 35.970 48.590 ;
        RECT 37.460 48.950 37.840 49.000 ;
        RECT 37.460 48.590 38.790 48.950 ;
        RECT 37.460 48.540 37.840 48.590 ;
      LAYER mcon ;
        RECT 18.855 49.980 19.155 50.280 ;
        RECT 33.230 49.980 33.530 50.280 ;
        RECT 27.970 48.620 28.270 48.920 ;
        RECT 28.460 48.620 28.760 48.920 ;
        RECT 28.950 48.620 29.250 48.920 ;
        RECT 34.640 48.620 34.940 48.920 ;
        RECT 35.130 48.620 35.430 48.920 ;
        RECT 35.620 48.620 35.920 48.920 ;
        RECT 37.510 48.620 37.810 48.920 ;
        RECT 38.000 48.620 38.300 48.920 ;
        RECT 38.490 48.620 38.790 48.920 ;
      LAYER met1 ;
        RECT 18.795 49.950 35.550 50.310 ;
        RECT 28.460 48.950 28.820 49.950 ;
        RECT 35.190 48.950 35.550 49.950 ;
        RECT 27.910 48.590 29.410 48.950 ;
        RECT 34.580 48.590 38.850 48.950 ;
      LAYER via ;
        RECT 27.110 49.950 27.470 50.310 ;
      LAYER met2 ;
        RECT 27.080 49.950 27.500 57.500 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 36.565 42.500 36.865 55.090 ;
        RECT 46.630 48.950 47.010 49.000 ;
        RECT 45.680 48.590 47.010 48.950 ;
        RECT 46.630 48.540 47.010 48.590 ;
        RECT 50.940 42.500 51.240 55.090 ;
        RECT 53.300 48.950 53.680 49.000 ;
        RECT 52.350 48.590 53.680 48.950 ;
        RECT 53.300 48.540 53.680 48.590 ;
        RECT 55.170 48.950 55.550 49.000 ;
        RECT 55.170 48.590 56.500 48.950 ;
        RECT 55.170 48.540 55.550 48.590 ;
      LAYER mcon ;
        RECT 36.565 49.980 36.865 50.280 ;
        RECT 50.940 49.980 51.240 50.280 ;
        RECT 45.680 48.620 45.980 48.920 ;
        RECT 46.170 48.620 46.470 48.920 ;
        RECT 46.660 48.620 46.960 48.920 ;
        RECT 52.350 48.620 52.650 48.920 ;
        RECT 52.840 48.620 53.140 48.920 ;
        RECT 53.330 48.620 53.630 48.920 ;
        RECT 55.220 48.620 55.520 48.920 ;
        RECT 55.710 48.620 56.010 48.920 ;
        RECT 56.200 48.620 56.500 48.920 ;
      LAYER met1 ;
        RECT 36.505 49.950 53.260 50.310 ;
        RECT 46.170 48.950 46.530 49.950 ;
        RECT 52.900 48.950 53.260 49.950 ;
        RECT 45.620 48.590 47.120 48.950 ;
        RECT 52.290 48.590 56.560 48.950 ;
      LAYER via ;
        RECT 51.480 49.950 51.840 50.310 ;
      LAYER met2 ;
        RECT 51.450 49.950 51.870 57.500 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 54.275 42.500 54.575 55.090 ;
        RECT 64.340 48.950 64.720 49.000 ;
        RECT 63.390 48.590 64.720 48.950 ;
        RECT 64.340 48.540 64.720 48.590 ;
        RECT 68.650 42.500 68.950 55.090 ;
        RECT 71.010 48.950 71.390 49.000 ;
        RECT 70.060 48.590 71.390 48.950 ;
        RECT 71.010 48.540 71.390 48.590 ;
        RECT 72.880 48.950 73.260 49.000 ;
        RECT 72.880 48.590 74.210 48.950 ;
        RECT 72.880 48.540 73.260 48.590 ;
      LAYER mcon ;
        RECT 54.275 49.980 54.575 50.280 ;
        RECT 68.650 49.980 68.950 50.280 ;
        RECT 63.390 48.620 63.690 48.920 ;
        RECT 63.880 48.620 64.180 48.920 ;
        RECT 64.370 48.620 64.670 48.920 ;
        RECT 70.060 48.620 70.360 48.920 ;
        RECT 70.550 48.620 70.850 48.920 ;
        RECT 71.040 48.620 71.340 48.920 ;
        RECT 72.930 48.620 73.230 48.920 ;
        RECT 73.420 48.620 73.720 48.920 ;
        RECT 73.910 48.620 74.210 48.920 ;
      LAYER met1 ;
        RECT 54.215 49.950 70.970 50.310 ;
        RECT 63.880 48.950 64.240 49.950 ;
        RECT 70.610 48.950 70.970 49.950 ;
        RECT 63.330 48.590 64.830 48.950 ;
        RECT 70.000 48.590 74.270 48.950 ;
      LAYER via ;
        RECT 68.270 49.950 68.630 50.310 ;
      LAYER met2 ;
        RECT 68.240 49.950 68.660 57.500 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 71.985 42.500 72.285 55.090 ;
        RECT 82.050 48.950 82.430 49.000 ;
        RECT 81.100 48.590 82.430 48.950 ;
        RECT 82.050 48.540 82.430 48.590 ;
        RECT 86.360 42.500 86.660 55.090 ;
        RECT 88.720 48.950 89.100 49.000 ;
        RECT 87.770 48.590 89.100 48.950 ;
        RECT 88.720 48.540 89.100 48.590 ;
        RECT 90.590 48.950 90.970 49.000 ;
        RECT 90.590 48.590 91.920 48.950 ;
        RECT 90.590 48.540 90.970 48.590 ;
      LAYER mcon ;
        RECT 71.985 49.980 72.285 50.280 ;
        RECT 86.360 49.980 86.660 50.280 ;
        RECT 81.100 48.620 81.400 48.920 ;
        RECT 81.590 48.620 81.890 48.920 ;
        RECT 82.080 48.620 82.380 48.920 ;
        RECT 87.770 48.620 88.070 48.920 ;
        RECT 88.260 48.620 88.560 48.920 ;
        RECT 88.750 48.620 89.050 48.920 ;
        RECT 90.640 48.620 90.940 48.920 ;
        RECT 91.130 48.620 91.430 48.920 ;
        RECT 91.620 48.620 91.920 48.920 ;
      LAYER met1 ;
        RECT 71.925 49.950 88.680 50.310 ;
        RECT 81.590 48.950 81.950 49.950 ;
        RECT 88.320 48.950 88.680 49.950 ;
        RECT 81.040 48.590 82.540 48.950 ;
        RECT 87.710 48.590 91.980 48.950 ;
      LAYER via ;
        RECT 83.570 49.950 83.930 50.310 ;
      LAYER met2 ;
        RECT 83.540 49.950 83.960 57.500 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 89.695 42.500 89.995 55.090 ;
        RECT 99.760 48.950 100.140 49.000 ;
        RECT 98.810 48.590 100.140 48.950 ;
        RECT 99.760 48.540 100.140 48.590 ;
        RECT 104.070 42.500 104.370 55.090 ;
        RECT 110.130 33.250 110.510 33.300 ;
        RECT 109.180 32.890 110.510 33.250 ;
        RECT 110.130 32.840 110.510 32.890 ;
        RECT 112.000 33.250 112.380 33.300 ;
        RECT 112.000 32.890 113.330 33.250 ;
        RECT 112.000 32.840 112.380 32.890 ;
      LAYER mcon ;
        RECT 89.695 49.980 89.995 50.280 ;
        RECT 104.070 49.980 104.370 50.280 ;
        RECT 98.810 48.620 99.110 48.920 ;
        RECT 99.300 48.620 99.600 48.920 ;
        RECT 99.790 48.620 100.090 48.920 ;
        RECT 109.180 32.920 109.480 33.220 ;
        RECT 109.670 32.920 109.970 33.220 ;
        RECT 110.160 32.920 110.460 33.220 ;
        RECT 112.050 32.920 112.350 33.220 ;
        RECT 112.540 32.920 112.840 33.220 ;
        RECT 113.030 32.920 113.330 33.220 ;
      LAYER met1 ;
        RECT 89.635 49.950 107.720 50.310 ;
        RECT 99.300 48.950 99.660 49.950 ;
        RECT 98.750 48.590 100.250 48.950 ;
        RECT 107.360 43.360 107.720 49.950 ;
        RECT 107.360 43.000 116.860 43.360 ;
        RECT 109.120 32.890 113.390 33.250 ;
        RECT 112.420 31.890 112.780 32.890 ;
        RECT 116.500 31.890 116.860 43.000 ;
        RECT 112.420 31.530 116.860 31.890 ;
      LAYER via ;
        RECT 106.000 49.950 106.360 50.310 ;
      LAYER met2 ;
        RECT 105.970 49.950 106.390 57.500 ;
    END
  END p[10]
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 6.775 50.300 7.235 50.525 ;
        RECT -0.400 50.000 7.235 50.300 ;
        RECT 6.775 49.795 7.235 50.000 ;
      LAYER mcon ;
        RECT -0.380 50.020 -0.120 50.280 ;
      LAYER met1 ;
        RECT -0.450 49.950 -0.050 50.350 ;
    END
  END enb
  PIN input_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 115.015 44.500 116.000 45.500 ;
        RECT 115.015 43.500 115.380 44.500 ;
      LAYER mcon ;
        RECT 115.105 45.100 115.405 45.400 ;
        RECT 115.595 45.100 115.895 45.400 ;
        RECT 115.105 44.600 115.405 44.900 ;
        RECT 115.595 44.600 115.895 44.900 ;
      LAYER met1 ;
        RECT 115.015 44.500 116.000 45.500 ;
        RECT 122.630 45.030 123.070 45.470 ;
      LAYER via ;
        RECT 115.085 45.080 115.425 45.420 ;
        RECT 115.575 45.080 115.915 45.420 ;
        RECT 122.660 45.060 123.040 45.440 ;
        RECT 115.085 44.580 115.425 44.920 ;
        RECT 115.575 44.580 115.915 44.920 ;
      LAYER met2 ;
        RECT 115.015 45.000 123.100 45.500 ;
        RECT 115.015 44.500 116.000 45.000 ;
      LAYER via2 ;
        RECT 122.650 45.050 123.050 45.450 ;
      LAYER met3 ;
        RECT 122.570 44.970 123.130 45.530 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.500 50.105 9.180 51.950 ;
        RECT 10.495 50.105 12.255 51.950 ;
        RECT 15.980 48.965 105.050 55.840 ;
        RECT 27.020 48.960 34.210 48.965 ;
        RECT 44.730 48.960 51.920 48.965 ;
        RECT 62.440 48.960 69.630 48.965 ;
        RECT 80.150 48.960 87.340 48.965 ;
        RECT 97.860 48.960 105.050 48.965 ;
        RECT 7.500 32.875 14.690 32.880 ;
        RECT 25.210 32.875 32.400 32.880 ;
        RECT 42.920 32.875 50.110 32.880 ;
        RECT 60.630 32.875 67.820 32.880 ;
        RECT 78.340 32.875 85.530 32.880 ;
        RECT 96.050 32.875 103.240 32.880 ;
        RECT 7.500 26.000 114.280 32.875 ;
      LAYER li1 ;
        RECT 16.160 55.660 18.050 55.690 ;
        RECT 19.840 55.660 23.690 55.690 ;
        RECT 25.350 55.660 29.200 55.690 ;
        RECT 31.040 55.660 32.440 55.690 ;
        RECT 33.870 55.660 35.760 55.690 ;
        RECT 37.550 55.660 41.400 55.690 ;
        RECT 43.060 55.660 46.910 55.690 ;
        RECT 48.750 55.660 50.150 55.690 ;
        RECT 51.580 55.660 53.470 55.690 ;
        RECT 55.260 55.660 59.110 55.690 ;
        RECT 60.770 55.660 64.620 55.690 ;
        RECT 66.460 55.660 67.860 55.690 ;
        RECT 69.290 55.660 71.180 55.690 ;
        RECT 72.970 55.660 76.820 55.690 ;
        RECT 78.480 55.660 82.330 55.690 ;
        RECT 84.170 55.660 85.570 55.690 ;
        RECT 87.000 55.660 88.890 55.690 ;
        RECT 90.680 55.660 94.530 55.690 ;
        RECT 96.190 55.660 100.040 55.690 ;
        RECT 101.880 55.660 103.280 55.690 ;
        RECT 16.160 55.490 104.870 55.660 ;
        RECT 16.160 55.330 18.050 55.490 ;
        RECT 19.840 55.330 23.690 55.490 ;
        RECT 25.350 55.330 29.200 55.490 ;
        RECT 31.040 55.330 32.440 55.490 ;
        RECT 33.870 55.330 35.760 55.490 ;
        RECT 37.550 55.330 41.400 55.490 ;
        RECT 43.060 55.330 46.910 55.490 ;
        RECT 48.750 55.330 50.150 55.490 ;
        RECT 51.580 55.330 53.470 55.490 ;
        RECT 55.260 55.330 59.110 55.490 ;
        RECT 60.770 55.330 64.620 55.490 ;
        RECT 66.460 55.330 67.860 55.490 ;
        RECT 69.290 55.330 71.180 55.490 ;
        RECT 72.970 55.330 76.820 55.490 ;
        RECT 78.480 55.330 82.330 55.490 ;
        RECT 84.170 55.330 85.570 55.490 ;
        RECT 87.000 55.330 88.890 55.490 ;
        RECT 90.680 55.330 94.530 55.490 ;
        RECT 96.190 55.330 100.040 55.490 ;
        RECT 101.880 55.330 103.280 55.490 ;
        RECT 6.690 51.605 7.690 51.770 ;
        RECT 10.685 51.605 11.685 51.770 ;
        RECT 6.690 51.435 8.990 51.605 ;
        RECT 10.685 51.435 12.065 51.605 ;
        RECT 7.205 51.035 8.140 51.435 ;
        RECT 10.960 50.710 11.290 51.435 ;
        RECT 16.160 50.460 16.330 55.330 ;
        RECT 16.670 50.040 16.960 55.330 ;
        RECT 21.050 50.040 21.340 55.330 ;
        RECT 21.680 50.460 21.850 55.330 ;
        RECT 22.190 50.040 22.480 55.330 ;
        RECT 26.570 50.040 26.860 55.330 ;
        RECT 27.200 50.460 27.370 55.330 ;
        RECT 27.710 50.030 28.000 55.330 ;
        RECT 31.040 50.030 31.330 55.330 ;
        RECT 33.870 50.460 34.040 55.330 ;
        RECT 34.380 50.040 34.670 55.330 ;
        RECT 38.760 50.040 39.050 55.330 ;
        RECT 39.390 50.460 39.560 55.330 ;
        RECT 39.900 50.040 40.190 55.330 ;
        RECT 44.280 50.040 44.570 55.330 ;
        RECT 44.910 50.460 45.080 55.330 ;
        RECT 45.420 50.030 45.710 55.330 ;
        RECT 48.750 50.030 49.040 55.330 ;
        RECT 51.580 50.460 51.750 55.330 ;
        RECT 52.090 50.040 52.380 55.330 ;
        RECT 56.470 50.040 56.760 55.330 ;
        RECT 57.100 50.460 57.270 55.330 ;
        RECT 57.610 50.040 57.900 55.330 ;
        RECT 61.990 50.040 62.280 55.330 ;
        RECT 62.620 50.460 62.790 55.330 ;
        RECT 63.130 50.030 63.420 55.330 ;
        RECT 66.460 50.030 66.750 55.330 ;
        RECT 69.290 50.460 69.460 55.330 ;
        RECT 69.800 50.040 70.090 55.330 ;
        RECT 74.180 50.040 74.470 55.330 ;
        RECT 74.810 50.460 74.980 55.330 ;
        RECT 75.320 50.040 75.610 55.330 ;
        RECT 79.700 50.040 79.990 55.330 ;
        RECT 80.330 50.460 80.500 55.330 ;
        RECT 80.840 50.030 81.130 55.330 ;
        RECT 84.170 50.030 84.460 55.330 ;
        RECT 87.000 50.460 87.170 55.330 ;
        RECT 87.510 50.040 87.800 55.330 ;
        RECT 91.890 50.040 92.180 55.330 ;
        RECT 92.520 50.460 92.690 55.330 ;
        RECT 93.030 50.040 93.320 55.330 ;
        RECT 97.410 50.040 97.700 55.330 ;
        RECT 98.040 50.460 98.210 55.330 ;
        RECT 98.550 50.030 98.840 55.330 ;
        RECT 101.880 50.030 102.170 55.330 ;
        RECT 10.380 26.510 10.670 31.810 ;
        RECT 13.710 26.510 14.000 31.810 ;
        RECT 14.340 26.510 14.510 31.380 ;
        RECT 14.850 26.510 15.140 31.800 ;
        RECT 19.230 26.510 19.520 31.800 ;
        RECT 19.860 26.510 20.030 31.380 ;
        RECT 20.370 26.510 20.660 31.800 ;
        RECT 24.750 26.510 25.040 31.800 ;
        RECT 25.380 26.510 25.550 31.380 ;
        RECT 28.090 26.510 28.380 31.810 ;
        RECT 31.420 26.510 31.710 31.810 ;
        RECT 32.050 26.510 32.220 31.380 ;
        RECT 32.560 26.510 32.850 31.800 ;
        RECT 36.940 26.510 37.230 31.800 ;
        RECT 37.570 26.510 37.740 31.380 ;
        RECT 38.080 26.510 38.370 31.800 ;
        RECT 42.460 26.510 42.750 31.800 ;
        RECT 43.090 26.510 43.260 31.380 ;
        RECT 45.800 26.510 46.090 31.810 ;
        RECT 49.130 26.510 49.420 31.810 ;
        RECT 49.760 26.510 49.930 31.380 ;
        RECT 50.270 26.510 50.560 31.800 ;
        RECT 54.650 26.510 54.940 31.800 ;
        RECT 55.280 26.510 55.450 31.380 ;
        RECT 55.790 26.510 56.080 31.800 ;
        RECT 60.170 26.510 60.460 31.800 ;
        RECT 60.800 26.510 60.970 31.380 ;
        RECT 63.510 26.510 63.800 31.810 ;
        RECT 66.840 26.510 67.130 31.810 ;
        RECT 67.470 26.510 67.640 31.380 ;
        RECT 67.980 26.510 68.270 31.800 ;
        RECT 72.360 26.510 72.650 31.800 ;
        RECT 72.990 26.510 73.160 31.380 ;
        RECT 73.500 26.510 73.790 31.800 ;
        RECT 77.880 26.510 78.170 31.800 ;
        RECT 78.510 26.510 78.680 31.380 ;
        RECT 81.220 26.510 81.510 31.810 ;
        RECT 84.550 26.510 84.840 31.810 ;
        RECT 85.180 26.510 85.350 31.380 ;
        RECT 85.690 26.510 85.980 31.800 ;
        RECT 90.070 26.510 90.360 31.800 ;
        RECT 90.700 26.510 90.870 31.380 ;
        RECT 91.210 26.510 91.500 31.800 ;
        RECT 95.590 26.510 95.880 31.800 ;
        RECT 96.220 26.510 96.390 31.380 ;
        RECT 98.930 26.510 99.220 31.810 ;
        RECT 102.260 26.510 102.550 31.810 ;
        RECT 102.890 26.510 103.060 31.380 ;
        RECT 103.400 26.510 103.690 31.800 ;
        RECT 107.780 26.510 108.070 31.800 ;
        RECT 108.410 26.510 108.580 31.380 ;
        RECT 108.920 26.510 109.210 31.800 ;
        RECT 113.300 26.510 113.590 31.800 ;
        RECT 113.930 26.510 114.100 31.380 ;
        RECT 9.270 26.350 10.670 26.510 ;
        RECT 12.510 26.350 16.360 26.510 ;
        RECT 18.020 26.350 21.870 26.510 ;
        RECT 23.660 26.350 25.550 26.510 ;
        RECT 26.980 26.350 28.380 26.510 ;
        RECT 30.220 26.350 34.070 26.510 ;
        RECT 35.730 26.350 39.580 26.510 ;
        RECT 41.370 26.350 43.260 26.510 ;
        RECT 44.690 26.350 46.090 26.510 ;
        RECT 47.930 26.350 51.780 26.510 ;
        RECT 53.440 26.350 57.290 26.510 ;
        RECT 59.080 26.350 60.970 26.510 ;
        RECT 62.400 26.350 63.800 26.510 ;
        RECT 65.640 26.350 69.490 26.510 ;
        RECT 71.150 26.350 75.000 26.510 ;
        RECT 76.790 26.350 78.680 26.510 ;
        RECT 80.110 26.350 81.510 26.510 ;
        RECT 83.350 26.350 87.200 26.510 ;
        RECT 88.860 26.350 92.710 26.510 ;
        RECT 94.500 26.350 96.390 26.510 ;
        RECT 97.820 26.350 99.220 26.510 ;
        RECT 101.060 26.350 104.910 26.510 ;
        RECT 106.570 26.350 110.420 26.510 ;
        RECT 112.210 26.350 114.100 26.510 ;
        RECT 7.680 26.180 114.100 26.350 ;
        RECT 9.270 26.150 10.670 26.180 ;
        RECT 12.510 26.150 16.360 26.180 ;
        RECT 18.020 26.150 21.870 26.180 ;
        RECT 23.660 26.150 25.550 26.180 ;
        RECT 26.980 26.150 28.380 26.180 ;
        RECT 30.220 26.150 34.070 26.180 ;
        RECT 35.730 26.150 39.580 26.180 ;
        RECT 41.370 26.150 43.260 26.180 ;
        RECT 44.690 26.150 46.090 26.180 ;
        RECT 47.930 26.150 51.780 26.180 ;
        RECT 53.440 26.150 57.290 26.180 ;
        RECT 59.080 26.150 60.970 26.180 ;
        RECT 62.400 26.150 63.800 26.180 ;
        RECT 65.640 26.150 69.490 26.180 ;
        RECT 71.150 26.150 75.000 26.180 ;
        RECT 76.790 26.150 78.680 26.180 ;
        RECT 80.110 26.150 81.510 26.180 ;
        RECT 83.350 26.150 87.200 26.180 ;
        RECT 88.860 26.150 92.710 26.180 ;
        RECT 94.500 26.150 96.390 26.180 ;
        RECT 97.820 26.150 99.220 26.180 ;
        RECT 101.060 26.150 104.910 26.180 ;
        RECT 106.570 26.150 110.420 26.180 ;
        RECT 112.210 26.150 114.100 26.180 ;
      LAYER mcon ;
        RECT 16.220 55.360 16.520 55.660 ;
        RECT 16.710 55.360 17.010 55.660 ;
        RECT 17.200 55.360 17.500 55.660 ;
        RECT 17.690 55.360 17.990 55.660 ;
        RECT 19.900 55.360 20.200 55.660 ;
        RECT 20.390 55.360 20.690 55.660 ;
        RECT 20.880 55.360 21.180 55.660 ;
        RECT 21.370 55.360 21.670 55.660 ;
        RECT 21.860 55.360 22.160 55.660 ;
        RECT 22.350 55.360 22.650 55.660 ;
        RECT 22.840 55.360 23.140 55.660 ;
        RECT 23.330 55.360 23.630 55.660 ;
        RECT 25.410 55.360 25.710 55.660 ;
        RECT 25.900 55.360 26.200 55.660 ;
        RECT 26.390 55.360 26.690 55.660 ;
        RECT 26.880 55.360 27.180 55.660 ;
        RECT 27.370 55.360 27.670 55.660 ;
        RECT 27.860 55.360 28.160 55.660 ;
        RECT 28.350 55.360 28.650 55.660 ;
        RECT 28.840 55.360 29.140 55.660 ;
        RECT 31.100 55.360 31.400 55.660 ;
        RECT 31.590 55.360 31.890 55.660 ;
        RECT 32.080 55.360 32.380 55.660 ;
        RECT 33.930 55.360 34.230 55.660 ;
        RECT 34.420 55.360 34.720 55.660 ;
        RECT 34.910 55.360 35.210 55.660 ;
        RECT 35.400 55.360 35.700 55.660 ;
        RECT 37.610 55.360 37.910 55.660 ;
        RECT 38.100 55.360 38.400 55.660 ;
        RECT 38.590 55.360 38.890 55.660 ;
        RECT 39.080 55.360 39.380 55.660 ;
        RECT 39.570 55.360 39.870 55.660 ;
        RECT 40.060 55.360 40.360 55.660 ;
        RECT 40.550 55.360 40.850 55.660 ;
        RECT 41.040 55.360 41.340 55.660 ;
        RECT 43.120 55.360 43.420 55.660 ;
        RECT 43.610 55.360 43.910 55.660 ;
        RECT 44.100 55.360 44.400 55.660 ;
        RECT 44.590 55.360 44.890 55.660 ;
        RECT 45.080 55.360 45.380 55.660 ;
        RECT 45.570 55.360 45.870 55.660 ;
        RECT 46.060 55.360 46.360 55.660 ;
        RECT 46.550 55.360 46.850 55.660 ;
        RECT 48.810 55.360 49.110 55.660 ;
        RECT 49.300 55.360 49.600 55.660 ;
        RECT 49.790 55.360 50.090 55.660 ;
        RECT 51.640 55.360 51.940 55.660 ;
        RECT 52.130 55.360 52.430 55.660 ;
        RECT 52.620 55.360 52.920 55.660 ;
        RECT 53.110 55.360 53.410 55.660 ;
        RECT 55.320 55.360 55.620 55.660 ;
        RECT 55.810 55.360 56.110 55.660 ;
        RECT 56.300 55.360 56.600 55.660 ;
        RECT 56.790 55.360 57.090 55.660 ;
        RECT 57.280 55.360 57.580 55.660 ;
        RECT 57.770 55.360 58.070 55.660 ;
        RECT 58.260 55.360 58.560 55.660 ;
        RECT 58.750 55.360 59.050 55.660 ;
        RECT 60.830 55.360 61.130 55.660 ;
        RECT 61.320 55.360 61.620 55.660 ;
        RECT 61.810 55.360 62.110 55.660 ;
        RECT 62.300 55.360 62.600 55.660 ;
        RECT 62.790 55.360 63.090 55.660 ;
        RECT 63.280 55.360 63.580 55.660 ;
        RECT 63.770 55.360 64.070 55.660 ;
        RECT 64.260 55.360 64.560 55.660 ;
        RECT 66.520 55.360 66.820 55.660 ;
        RECT 67.010 55.360 67.310 55.660 ;
        RECT 67.500 55.360 67.800 55.660 ;
        RECT 69.350 55.360 69.650 55.660 ;
        RECT 69.840 55.360 70.140 55.660 ;
        RECT 70.330 55.360 70.630 55.660 ;
        RECT 70.820 55.360 71.120 55.660 ;
        RECT 73.030 55.360 73.330 55.660 ;
        RECT 73.520 55.360 73.820 55.660 ;
        RECT 74.010 55.360 74.310 55.660 ;
        RECT 74.500 55.360 74.800 55.660 ;
        RECT 74.990 55.360 75.290 55.660 ;
        RECT 75.480 55.360 75.780 55.660 ;
        RECT 75.970 55.360 76.270 55.660 ;
        RECT 76.460 55.360 76.760 55.660 ;
        RECT 78.540 55.360 78.840 55.660 ;
        RECT 79.030 55.360 79.330 55.660 ;
        RECT 79.520 55.360 79.820 55.660 ;
        RECT 80.010 55.360 80.310 55.660 ;
        RECT 80.500 55.360 80.800 55.660 ;
        RECT 80.990 55.360 81.290 55.660 ;
        RECT 81.480 55.360 81.780 55.660 ;
        RECT 81.970 55.360 82.270 55.660 ;
        RECT 84.230 55.360 84.530 55.660 ;
        RECT 84.720 55.360 85.020 55.660 ;
        RECT 85.210 55.360 85.510 55.660 ;
        RECT 87.060 55.360 87.360 55.660 ;
        RECT 87.550 55.360 87.850 55.660 ;
        RECT 88.040 55.360 88.340 55.660 ;
        RECT 88.530 55.360 88.830 55.660 ;
        RECT 90.740 55.360 91.040 55.660 ;
        RECT 91.230 55.360 91.530 55.660 ;
        RECT 91.720 55.360 92.020 55.660 ;
        RECT 92.210 55.360 92.510 55.660 ;
        RECT 92.700 55.360 93.000 55.660 ;
        RECT 93.190 55.360 93.490 55.660 ;
        RECT 93.680 55.360 93.980 55.660 ;
        RECT 94.170 55.360 94.470 55.660 ;
        RECT 96.250 55.360 96.550 55.660 ;
        RECT 96.740 55.360 97.040 55.660 ;
        RECT 97.230 55.360 97.530 55.660 ;
        RECT 97.720 55.360 98.020 55.660 ;
        RECT 98.210 55.360 98.510 55.660 ;
        RECT 98.700 55.360 99.000 55.660 ;
        RECT 99.190 55.360 99.490 55.660 ;
        RECT 99.680 55.360 99.980 55.660 ;
        RECT 101.940 55.360 102.240 55.660 ;
        RECT 102.430 55.360 102.730 55.660 ;
        RECT 102.920 55.360 103.220 55.660 ;
        RECT 6.835 51.435 7.005 51.605 ;
        RECT 7.295 51.435 7.465 51.605 ;
        RECT 7.755 51.435 7.925 51.605 ;
        RECT 8.215 51.435 8.385 51.605 ;
        RECT 8.675 51.435 8.845 51.605 ;
        RECT 10.830 51.435 11.000 51.605 ;
        RECT 11.290 51.435 11.460 51.605 ;
        RECT 11.750 51.435 11.920 51.605 ;
        RECT 9.330 26.180 9.630 26.480 ;
        RECT 9.820 26.180 10.120 26.480 ;
        RECT 10.310 26.180 10.610 26.480 ;
        RECT 12.570 26.180 12.870 26.480 ;
        RECT 13.060 26.180 13.360 26.480 ;
        RECT 13.550 26.180 13.850 26.480 ;
        RECT 14.040 26.180 14.340 26.480 ;
        RECT 14.530 26.180 14.830 26.480 ;
        RECT 15.020 26.180 15.320 26.480 ;
        RECT 15.510 26.180 15.810 26.480 ;
        RECT 16.000 26.180 16.300 26.480 ;
        RECT 18.080 26.180 18.380 26.480 ;
        RECT 18.570 26.180 18.870 26.480 ;
        RECT 19.060 26.180 19.360 26.480 ;
        RECT 19.550 26.180 19.850 26.480 ;
        RECT 20.040 26.180 20.340 26.480 ;
        RECT 20.530 26.180 20.830 26.480 ;
        RECT 21.020 26.180 21.320 26.480 ;
        RECT 21.510 26.180 21.810 26.480 ;
        RECT 23.720 26.180 24.020 26.480 ;
        RECT 24.210 26.180 24.510 26.480 ;
        RECT 24.700 26.180 25.000 26.480 ;
        RECT 25.190 26.180 25.490 26.480 ;
        RECT 27.040 26.180 27.340 26.480 ;
        RECT 27.530 26.180 27.830 26.480 ;
        RECT 28.020 26.180 28.320 26.480 ;
        RECT 30.280 26.180 30.580 26.480 ;
        RECT 30.770 26.180 31.070 26.480 ;
        RECT 31.260 26.180 31.560 26.480 ;
        RECT 31.750 26.180 32.050 26.480 ;
        RECT 32.240 26.180 32.540 26.480 ;
        RECT 32.730 26.180 33.030 26.480 ;
        RECT 33.220 26.180 33.520 26.480 ;
        RECT 33.710 26.180 34.010 26.480 ;
        RECT 35.790 26.180 36.090 26.480 ;
        RECT 36.280 26.180 36.580 26.480 ;
        RECT 36.770 26.180 37.070 26.480 ;
        RECT 37.260 26.180 37.560 26.480 ;
        RECT 37.750 26.180 38.050 26.480 ;
        RECT 38.240 26.180 38.540 26.480 ;
        RECT 38.730 26.180 39.030 26.480 ;
        RECT 39.220 26.180 39.520 26.480 ;
        RECT 41.430 26.180 41.730 26.480 ;
        RECT 41.920 26.180 42.220 26.480 ;
        RECT 42.410 26.180 42.710 26.480 ;
        RECT 42.900 26.180 43.200 26.480 ;
        RECT 44.750 26.180 45.050 26.480 ;
        RECT 45.240 26.180 45.540 26.480 ;
        RECT 45.730 26.180 46.030 26.480 ;
        RECT 47.990 26.180 48.290 26.480 ;
        RECT 48.480 26.180 48.780 26.480 ;
        RECT 48.970 26.180 49.270 26.480 ;
        RECT 49.460 26.180 49.760 26.480 ;
        RECT 49.950 26.180 50.250 26.480 ;
        RECT 50.440 26.180 50.740 26.480 ;
        RECT 50.930 26.180 51.230 26.480 ;
        RECT 51.420 26.180 51.720 26.480 ;
        RECT 53.500 26.180 53.800 26.480 ;
        RECT 53.990 26.180 54.290 26.480 ;
        RECT 54.480 26.180 54.780 26.480 ;
        RECT 54.970 26.180 55.270 26.480 ;
        RECT 55.460 26.180 55.760 26.480 ;
        RECT 55.950 26.180 56.250 26.480 ;
        RECT 56.440 26.180 56.740 26.480 ;
        RECT 56.930 26.180 57.230 26.480 ;
        RECT 59.140 26.180 59.440 26.480 ;
        RECT 59.630 26.180 59.930 26.480 ;
        RECT 60.120 26.180 60.420 26.480 ;
        RECT 60.610 26.180 60.910 26.480 ;
        RECT 62.460 26.180 62.760 26.480 ;
        RECT 62.950 26.180 63.250 26.480 ;
        RECT 63.440 26.180 63.740 26.480 ;
        RECT 65.700 26.180 66.000 26.480 ;
        RECT 66.190 26.180 66.490 26.480 ;
        RECT 66.680 26.180 66.980 26.480 ;
        RECT 67.170 26.180 67.470 26.480 ;
        RECT 67.660 26.180 67.960 26.480 ;
        RECT 68.150 26.180 68.450 26.480 ;
        RECT 68.640 26.180 68.940 26.480 ;
        RECT 69.130 26.180 69.430 26.480 ;
        RECT 71.210 26.180 71.510 26.480 ;
        RECT 71.700 26.180 72.000 26.480 ;
        RECT 72.190 26.180 72.490 26.480 ;
        RECT 72.680 26.180 72.980 26.480 ;
        RECT 73.170 26.180 73.470 26.480 ;
        RECT 73.660 26.180 73.960 26.480 ;
        RECT 74.150 26.180 74.450 26.480 ;
        RECT 74.640 26.180 74.940 26.480 ;
        RECT 76.850 26.180 77.150 26.480 ;
        RECT 77.340 26.180 77.640 26.480 ;
        RECT 77.830 26.180 78.130 26.480 ;
        RECT 78.320 26.180 78.620 26.480 ;
        RECT 80.170 26.180 80.470 26.480 ;
        RECT 80.660 26.180 80.960 26.480 ;
        RECT 81.150 26.180 81.450 26.480 ;
        RECT 83.410 26.180 83.710 26.480 ;
        RECT 83.900 26.180 84.200 26.480 ;
        RECT 84.390 26.180 84.690 26.480 ;
        RECT 84.880 26.180 85.180 26.480 ;
        RECT 85.370 26.180 85.670 26.480 ;
        RECT 85.860 26.180 86.160 26.480 ;
        RECT 86.350 26.180 86.650 26.480 ;
        RECT 86.840 26.180 87.140 26.480 ;
        RECT 88.920 26.180 89.220 26.480 ;
        RECT 89.410 26.180 89.710 26.480 ;
        RECT 89.900 26.180 90.200 26.480 ;
        RECT 90.390 26.180 90.690 26.480 ;
        RECT 90.880 26.180 91.180 26.480 ;
        RECT 91.370 26.180 91.670 26.480 ;
        RECT 91.860 26.180 92.160 26.480 ;
        RECT 92.350 26.180 92.650 26.480 ;
        RECT 94.560 26.180 94.860 26.480 ;
        RECT 95.050 26.180 95.350 26.480 ;
        RECT 95.540 26.180 95.840 26.480 ;
        RECT 96.030 26.180 96.330 26.480 ;
        RECT 97.880 26.180 98.180 26.480 ;
        RECT 98.370 26.180 98.670 26.480 ;
        RECT 98.860 26.180 99.160 26.480 ;
        RECT 101.120 26.180 101.420 26.480 ;
        RECT 101.610 26.180 101.910 26.480 ;
        RECT 102.100 26.180 102.400 26.480 ;
        RECT 102.590 26.180 102.890 26.480 ;
        RECT 103.080 26.180 103.380 26.480 ;
        RECT 103.570 26.180 103.870 26.480 ;
        RECT 104.060 26.180 104.360 26.480 ;
        RECT 104.550 26.180 104.850 26.480 ;
        RECT 106.630 26.180 106.930 26.480 ;
        RECT 107.120 26.180 107.420 26.480 ;
        RECT 107.610 26.180 107.910 26.480 ;
        RECT 108.100 26.180 108.400 26.480 ;
        RECT 108.590 26.180 108.890 26.480 ;
        RECT 109.080 26.180 109.380 26.480 ;
        RECT 109.570 26.180 109.870 26.480 ;
        RECT 110.060 26.180 110.360 26.480 ;
        RECT 112.270 26.180 112.570 26.480 ;
        RECT 112.760 26.180 113.060 26.480 ;
        RECT 113.250 26.180 113.550 26.480 ;
        RECT 113.740 26.180 114.040 26.480 ;
      LAYER met1 ;
        RECT 15.900 55.270 105.050 55.750 ;
        RECT 0.000 51.280 12.065 51.760 ;
        RECT 7.500 26.090 114.280 26.570 ;
      LAYER via ;
        RECT 18.130 55.360 18.430 55.660 ;
        RECT 18.490 55.360 18.790 55.660 ;
        RECT 18.850 55.360 19.150 55.660 ;
        RECT 19.210 55.360 19.510 55.660 ;
        RECT 19.570 55.360 19.870 55.660 ;
        RECT 46.130 55.360 46.430 55.660 ;
        RECT 46.490 55.360 46.790 55.660 ;
        RECT 46.850 55.360 47.150 55.660 ;
        RECT 47.210 55.360 47.510 55.660 ;
        RECT 47.570 55.360 47.870 55.660 ;
        RECT 74.130 55.360 74.430 55.660 ;
        RECT 74.490 55.360 74.790 55.660 ;
        RECT 74.850 55.360 75.150 55.660 ;
        RECT 75.210 55.360 75.510 55.660 ;
        RECT 75.570 55.360 75.870 55.660 ;
        RECT 102.130 55.360 102.430 55.660 ;
        RECT 102.490 55.360 102.790 55.660 ;
        RECT 102.850 55.360 103.150 55.660 ;
        RECT 103.210 55.360 103.510 55.660 ;
        RECT 103.570 55.360 103.870 55.660 ;
        RECT 0.130 51.370 0.430 51.670 ;
        RECT 0.490 51.370 0.790 51.670 ;
        RECT 0.850 51.370 1.150 51.670 ;
        RECT 1.210 51.370 1.510 51.670 ;
        RECT 1.570 51.370 1.870 51.670 ;
        RECT 18.130 26.180 18.430 26.480 ;
        RECT 18.490 26.180 18.790 26.480 ;
        RECT 18.850 26.180 19.150 26.480 ;
        RECT 19.210 26.180 19.510 26.480 ;
        RECT 19.570 26.180 19.870 26.480 ;
        RECT 46.130 26.180 46.430 26.480 ;
        RECT 46.490 26.180 46.790 26.480 ;
        RECT 46.850 26.180 47.150 26.480 ;
        RECT 47.210 26.180 47.510 26.480 ;
        RECT 47.570 26.180 47.870 26.480 ;
        RECT 74.130 26.180 74.430 26.480 ;
        RECT 74.490 26.180 74.790 26.480 ;
        RECT 74.850 26.180 75.150 26.480 ;
        RECT 75.210 26.180 75.510 26.480 ;
        RECT 75.570 26.180 75.870 26.480 ;
        RECT 102.130 26.180 102.430 26.480 ;
        RECT 102.490 26.180 102.790 26.480 ;
        RECT 102.850 26.180 103.150 26.480 ;
        RECT 103.210 26.180 103.510 26.480 ;
        RECT 103.570 26.180 103.870 26.480 ;
      LAYER met2 ;
        RECT 18.000 55.270 20.000 55.750 ;
        RECT 46.000 55.270 48.000 55.750 ;
        RECT 74.000 55.270 76.000 55.750 ;
        RECT 102.000 55.270 104.000 55.750 ;
        RECT 0.000 51.280 2.000 51.760 ;
        RECT 18.000 26.090 20.000 26.570 ;
        RECT 46.000 26.090 48.000 26.570 ;
        RECT 74.000 26.090 76.000 26.570 ;
        RECT 102.000 26.090 104.000 26.570 ;
      LAYER via2 ;
        RECT 18.180 55.350 18.500 55.670 ;
        RECT 18.620 55.350 18.940 55.670 ;
        RECT 19.060 55.350 19.380 55.670 ;
        RECT 19.500 55.350 19.820 55.670 ;
        RECT 46.180 55.350 46.500 55.670 ;
        RECT 46.620 55.350 46.940 55.670 ;
        RECT 47.060 55.350 47.380 55.670 ;
        RECT 47.500 55.350 47.820 55.670 ;
        RECT 74.180 55.350 74.500 55.670 ;
        RECT 74.620 55.350 74.940 55.670 ;
        RECT 75.060 55.350 75.380 55.670 ;
        RECT 75.500 55.350 75.820 55.670 ;
        RECT 102.180 55.350 102.500 55.670 ;
        RECT 102.620 55.350 102.940 55.670 ;
        RECT 103.060 55.350 103.380 55.670 ;
        RECT 103.500 55.350 103.820 55.670 ;
        RECT 0.180 51.360 0.500 51.680 ;
        RECT 0.620 51.360 0.940 51.680 ;
        RECT 1.060 51.360 1.380 51.680 ;
        RECT 1.500 51.360 1.820 51.680 ;
        RECT 18.180 26.170 18.500 26.490 ;
        RECT 18.620 26.170 18.940 26.490 ;
        RECT 19.060 26.170 19.380 26.490 ;
        RECT 19.500 26.170 19.820 26.490 ;
        RECT 46.180 26.170 46.500 26.490 ;
        RECT 46.620 26.170 46.940 26.490 ;
        RECT 47.060 26.170 47.380 26.490 ;
        RECT 47.500 26.170 47.820 26.490 ;
        RECT 74.180 26.170 74.500 26.490 ;
        RECT 74.620 26.170 74.940 26.490 ;
        RECT 75.060 26.170 75.380 26.490 ;
        RECT 75.500 26.170 75.820 26.490 ;
        RECT 102.180 26.170 102.500 26.490 ;
        RECT 102.620 26.170 102.940 26.490 ;
        RECT 103.060 26.170 103.380 26.490 ;
        RECT 103.500 26.170 103.820 26.490 ;
      LAYER met3 ;
        RECT 0.000 91.000 122.000 93.000 ;
        RECT 18.000 55.270 20.000 55.750 ;
        RECT 46.000 55.270 48.000 55.750 ;
        RECT 74.000 55.270 76.000 55.750 ;
        RECT 102.000 55.270 104.000 55.750 ;
        RECT 0.000 51.280 2.000 51.760 ;
        RECT 18.000 26.090 20.000 26.570 ;
        RECT 46.000 26.090 48.000 26.570 ;
        RECT 74.000 26.090 76.000 26.570 ;
        RECT 102.000 26.090 104.000 26.570 ;
        RECT 0.000 -12.000 122.000 -10.000 ;
      LAYER via3 ;
        RECT 0.200 92.400 0.600 92.800 ;
        RECT 0.800 92.400 1.200 92.800 ;
        RECT 1.400 92.400 1.800 92.800 ;
        RECT 18.200 92.400 18.600 92.800 ;
        RECT 18.800 92.400 19.200 92.800 ;
        RECT 19.400 92.400 19.800 92.800 ;
        RECT 46.200 92.400 46.600 92.800 ;
        RECT 46.800 92.400 47.200 92.800 ;
        RECT 47.400 92.400 47.800 92.800 ;
        RECT 74.200 92.400 74.600 92.800 ;
        RECT 74.800 92.400 75.200 92.800 ;
        RECT 75.400 92.400 75.800 92.800 ;
        RECT 102.200 92.400 102.600 92.800 ;
        RECT 102.800 92.400 103.200 92.800 ;
        RECT 103.400 92.400 103.800 92.800 ;
        RECT 120.200 92.400 120.600 92.800 ;
        RECT 120.800 92.400 121.200 92.800 ;
        RECT 121.400 92.400 121.800 92.800 ;
        RECT 0.200 91.800 0.600 92.200 ;
        RECT 0.800 91.800 1.200 92.200 ;
        RECT 1.400 91.800 1.800 92.200 ;
        RECT 18.200 91.800 18.600 92.200 ;
        RECT 18.800 91.800 19.200 92.200 ;
        RECT 19.400 91.800 19.800 92.200 ;
        RECT 46.200 91.800 46.600 92.200 ;
        RECT 46.800 91.800 47.200 92.200 ;
        RECT 47.400 91.800 47.800 92.200 ;
        RECT 74.200 91.800 74.600 92.200 ;
        RECT 74.800 91.800 75.200 92.200 ;
        RECT 75.400 91.800 75.800 92.200 ;
        RECT 102.200 91.800 102.600 92.200 ;
        RECT 102.800 91.800 103.200 92.200 ;
        RECT 103.400 91.800 103.800 92.200 ;
        RECT 120.200 91.800 120.600 92.200 ;
        RECT 120.800 91.800 121.200 92.200 ;
        RECT 121.400 91.800 121.800 92.200 ;
        RECT 0.200 91.200 0.600 91.600 ;
        RECT 0.800 91.200 1.200 91.600 ;
        RECT 1.400 91.200 1.800 91.600 ;
        RECT 18.200 91.200 18.600 91.600 ;
        RECT 18.800 91.200 19.200 91.600 ;
        RECT 19.400 91.200 19.800 91.600 ;
        RECT 46.200 91.200 46.600 91.600 ;
        RECT 46.800 91.200 47.200 91.600 ;
        RECT 47.400 91.200 47.800 91.600 ;
        RECT 74.200 91.200 74.600 91.600 ;
        RECT 74.800 91.200 75.200 91.600 ;
        RECT 75.400 91.200 75.800 91.600 ;
        RECT 102.200 91.200 102.600 91.600 ;
        RECT 102.800 91.200 103.200 91.600 ;
        RECT 103.400 91.200 103.800 91.600 ;
        RECT 120.200 91.200 120.600 91.600 ;
        RECT 120.800 91.200 121.200 91.600 ;
        RECT 121.400 91.200 121.800 91.600 ;
        RECT 18.160 55.330 18.520 55.695 ;
        RECT 18.600 55.330 18.960 55.695 ;
        RECT 19.040 55.330 19.400 55.695 ;
        RECT 19.480 55.330 19.840 55.695 ;
        RECT 46.160 55.330 46.520 55.695 ;
        RECT 46.600 55.330 46.960 55.695 ;
        RECT 47.040 55.330 47.400 55.695 ;
        RECT 47.480 55.330 47.840 55.695 ;
        RECT 74.160 55.330 74.520 55.695 ;
        RECT 74.600 55.330 74.960 55.695 ;
        RECT 75.040 55.330 75.400 55.695 ;
        RECT 75.480 55.330 75.840 55.695 ;
        RECT 102.160 55.330 102.520 55.695 ;
        RECT 102.600 55.330 102.960 55.695 ;
        RECT 103.040 55.330 103.400 55.695 ;
        RECT 103.480 55.330 103.840 55.695 ;
        RECT 0.160 51.340 0.520 51.705 ;
        RECT 0.600 51.340 0.960 51.705 ;
        RECT 1.040 51.340 1.400 51.705 ;
        RECT 1.480 51.340 1.840 51.705 ;
        RECT 18.160 26.150 18.520 26.515 ;
        RECT 18.600 26.150 18.960 26.515 ;
        RECT 19.040 26.150 19.400 26.515 ;
        RECT 19.480 26.150 19.840 26.515 ;
        RECT 46.160 26.150 46.520 26.515 ;
        RECT 46.600 26.150 46.960 26.515 ;
        RECT 47.040 26.150 47.400 26.515 ;
        RECT 47.480 26.150 47.840 26.515 ;
        RECT 74.160 26.150 74.520 26.515 ;
        RECT 74.600 26.150 74.960 26.515 ;
        RECT 75.040 26.150 75.400 26.515 ;
        RECT 75.480 26.150 75.840 26.515 ;
        RECT 102.160 26.150 102.520 26.515 ;
        RECT 102.600 26.150 102.960 26.515 ;
        RECT 103.040 26.150 103.400 26.515 ;
        RECT 103.480 26.150 103.840 26.515 ;
        RECT 0.200 -10.600 0.600 -10.200 ;
        RECT 0.800 -10.600 1.200 -10.200 ;
        RECT 1.400 -10.600 1.800 -10.200 ;
        RECT 18.200 -10.600 18.600 -10.200 ;
        RECT 18.800 -10.600 19.200 -10.200 ;
        RECT 19.400 -10.600 19.800 -10.200 ;
        RECT 46.200 -10.600 46.600 -10.200 ;
        RECT 46.800 -10.600 47.200 -10.200 ;
        RECT 47.400 -10.600 47.800 -10.200 ;
        RECT 74.200 -10.600 74.600 -10.200 ;
        RECT 74.800 -10.600 75.200 -10.200 ;
        RECT 75.400 -10.600 75.800 -10.200 ;
        RECT 102.200 -10.600 102.600 -10.200 ;
        RECT 102.800 -10.600 103.200 -10.200 ;
        RECT 103.400 -10.600 103.800 -10.200 ;
        RECT 120.200 -10.600 120.600 -10.200 ;
        RECT 120.800 -10.600 121.200 -10.200 ;
        RECT 121.400 -10.600 121.800 -10.200 ;
        RECT 0.200 -11.200 0.600 -10.800 ;
        RECT 0.800 -11.200 1.200 -10.800 ;
        RECT 1.400 -11.200 1.800 -10.800 ;
        RECT 18.200 -11.200 18.600 -10.800 ;
        RECT 18.800 -11.200 19.200 -10.800 ;
        RECT 19.400 -11.200 19.800 -10.800 ;
        RECT 46.200 -11.200 46.600 -10.800 ;
        RECT 46.800 -11.200 47.200 -10.800 ;
        RECT 47.400 -11.200 47.800 -10.800 ;
        RECT 74.200 -11.200 74.600 -10.800 ;
        RECT 74.800 -11.200 75.200 -10.800 ;
        RECT 75.400 -11.200 75.800 -10.800 ;
        RECT 102.200 -11.200 102.600 -10.800 ;
        RECT 102.800 -11.200 103.200 -10.800 ;
        RECT 103.400 -11.200 103.800 -10.800 ;
        RECT 120.200 -11.200 120.600 -10.800 ;
        RECT 120.800 -11.200 121.200 -10.800 ;
        RECT 121.400 -11.200 121.800 -10.800 ;
        RECT 0.200 -11.800 0.600 -11.400 ;
        RECT 0.800 -11.800 1.200 -11.400 ;
        RECT 1.400 -11.800 1.800 -11.400 ;
        RECT 18.200 -11.800 18.600 -11.400 ;
        RECT 18.800 -11.800 19.200 -11.400 ;
        RECT 19.400 -11.800 19.800 -11.400 ;
        RECT 46.200 -11.800 46.600 -11.400 ;
        RECT 46.800 -11.800 47.200 -11.400 ;
        RECT 47.400 -11.800 47.800 -11.400 ;
        RECT 74.200 -11.800 74.600 -11.400 ;
        RECT 74.800 -11.800 75.200 -11.400 ;
        RECT 75.400 -11.800 75.800 -11.400 ;
        RECT 102.200 -11.800 102.600 -11.400 ;
        RECT 102.800 -11.800 103.200 -11.400 ;
        RECT 103.400 -11.800 103.800 -11.400 ;
        RECT 120.200 -11.800 120.600 -11.400 ;
        RECT 120.800 -11.800 121.200 -11.400 ;
        RECT 121.400 -11.800 121.800 -11.400 ;
      LAYER met4 ;
        RECT 0.000 -12.000 2.000 93.000 ;
        RECT 18.000 -12.000 20.000 93.000 ;
        RECT 46.000 -12.000 48.000 93.000 ;
        RECT 74.000 -12.000 76.000 93.000 ;
        RECT 102.000 -12.000 104.000 93.000 ;
        RECT 120.000 -12.000 122.000 93.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 15.000 56.700 106.000 57.000 ;
        RECT 7.205 48.885 8.140 49.285 ;
        RECT 11.460 48.885 11.800 49.545 ;
        RECT 6.690 48.715 8.990 48.885 ;
        RECT 10.685 48.715 12.065 48.885 ;
        RECT 15.000 41.070 15.300 56.700 ;
        RECT 105.700 41.070 106.000 56.700 ;
        RECT 108.500 50.015 110.500 50.380 ;
        RECT 6.700 40.770 115.825 41.070 ;
        RECT 6.700 25.200 7.000 40.770 ;
        RECT 115.500 40.700 115.825 40.770 ;
        RECT 115.500 25.200 115.800 40.700 ;
        RECT 6.700 24.900 115.800 25.200 ;
      LAYER mcon ;
        RECT 32.110 56.700 32.410 57.000 ;
        RECT 32.600 56.700 32.900 57.000 ;
        RECT 33.100 56.700 33.400 57.000 ;
        RECT 33.590 56.700 33.890 57.000 ;
        RECT 60.110 56.700 60.410 57.000 ;
        RECT 60.600 56.700 60.900 57.000 ;
        RECT 61.100 56.700 61.400 57.000 ;
        RECT 61.590 56.700 61.890 57.000 ;
        RECT 88.110 56.700 88.410 57.000 ;
        RECT 88.600 56.700 88.900 57.000 ;
        RECT 89.100 56.700 89.400 57.000 ;
        RECT 89.590 56.700 89.890 57.000 ;
        RECT 6.835 48.715 7.005 48.885 ;
        RECT 7.295 48.715 7.465 48.885 ;
        RECT 7.755 48.715 7.925 48.885 ;
        RECT 8.215 48.715 8.385 48.885 ;
        RECT 8.675 48.715 8.845 48.885 ;
        RECT 10.830 48.715 11.000 48.885 ;
        RECT 11.290 48.715 11.460 48.885 ;
        RECT 11.750 48.715 11.920 48.885 ;
        RECT 108.600 50.050 108.900 50.350 ;
        RECT 109.100 50.050 109.400 50.350 ;
        RECT 109.600 50.050 109.900 50.350 ;
        RECT 110.100 50.050 110.400 50.350 ;
        RECT 32.110 24.900 32.410 25.200 ;
        RECT 32.600 24.900 32.900 25.200 ;
        RECT 33.100 24.900 33.400 25.200 ;
        RECT 33.590 24.900 33.890 25.200 ;
        RECT 60.110 24.900 60.410 25.200 ;
        RECT 60.600 24.900 60.900 25.200 ;
        RECT 61.100 24.900 61.400 25.200 ;
        RECT 61.590 24.900 61.890 25.200 ;
      LAYER met1 ;
        RECT 32.080 56.610 33.920 57.090 ;
        RECT 60.080 56.610 61.920 57.090 ;
        RECT 88.080 56.610 89.920 57.090 ;
        RECT 116.130 50.380 117.870 50.440 ;
        RECT 108.500 50.020 118.000 50.380 ;
        RECT 108.500 50.015 110.505 50.020 ;
        RECT 116.130 49.960 117.870 50.020 ;
        RECT 4.000 48.560 12.065 49.040 ;
        RECT 32.080 24.810 33.920 25.290 ;
        RECT 60.080 24.810 61.920 25.290 ;
      LAYER via ;
        RECT 32.130 56.700 32.430 57.000 ;
        RECT 32.490 56.700 32.790 57.000 ;
        RECT 32.850 56.700 33.150 57.000 ;
        RECT 33.210 56.700 33.510 57.000 ;
        RECT 33.570 56.700 33.870 57.000 ;
        RECT 60.130 56.700 60.430 57.000 ;
        RECT 60.490 56.700 60.790 57.000 ;
        RECT 60.850 56.700 61.150 57.000 ;
        RECT 61.210 56.700 61.510 57.000 ;
        RECT 61.570 56.700 61.870 57.000 ;
        RECT 88.130 56.700 88.430 57.000 ;
        RECT 88.490 56.700 88.790 57.000 ;
        RECT 88.850 56.700 89.150 57.000 ;
        RECT 89.210 56.700 89.510 57.000 ;
        RECT 89.570 56.700 89.870 57.000 ;
        RECT 116.130 50.050 116.430 50.350 ;
        RECT 116.490 50.050 116.790 50.350 ;
        RECT 116.850 50.050 117.150 50.350 ;
        RECT 117.210 50.050 117.510 50.350 ;
        RECT 117.570 50.050 117.870 50.350 ;
        RECT 4.130 48.650 4.430 48.950 ;
        RECT 4.490 48.650 4.790 48.950 ;
        RECT 4.850 48.650 5.150 48.950 ;
        RECT 5.210 48.650 5.510 48.950 ;
        RECT 5.570 48.650 5.870 48.950 ;
        RECT 32.130 24.900 32.430 25.200 ;
        RECT 32.490 24.900 32.790 25.200 ;
        RECT 32.850 24.900 33.150 25.200 ;
        RECT 33.210 24.900 33.510 25.200 ;
        RECT 33.570 24.900 33.870 25.200 ;
        RECT 60.130 24.900 60.430 25.200 ;
        RECT 60.490 24.900 60.790 25.200 ;
        RECT 60.850 24.900 61.150 25.200 ;
        RECT 61.210 24.900 61.510 25.200 ;
        RECT 61.570 24.900 61.870 25.200 ;
      LAYER met2 ;
        RECT 32.000 56.610 34.000 57.090 ;
        RECT 60.000 56.610 62.000 57.090 ;
        RECT 88.000 56.610 90.000 57.090 ;
        RECT 116.000 49.960 118.000 50.440 ;
        RECT 4.000 48.560 6.000 49.040 ;
        RECT 32.000 24.810 34.000 25.290 ;
        RECT 60.000 24.810 62.000 25.290 ;
      LAYER via2 ;
        RECT 32.180 56.690 32.500 57.010 ;
        RECT 32.620 56.690 32.940 57.010 ;
        RECT 33.060 56.690 33.380 57.010 ;
        RECT 33.500 56.690 33.820 57.010 ;
        RECT 60.180 56.690 60.500 57.010 ;
        RECT 60.620 56.690 60.940 57.010 ;
        RECT 61.060 56.690 61.380 57.010 ;
        RECT 61.500 56.690 61.820 57.010 ;
        RECT 88.180 56.690 88.500 57.010 ;
        RECT 88.620 56.690 88.940 57.010 ;
        RECT 89.060 56.690 89.380 57.010 ;
        RECT 89.500 56.690 89.820 57.010 ;
        RECT 116.180 50.040 116.500 50.360 ;
        RECT 116.620 50.040 116.940 50.360 ;
        RECT 117.060 50.040 117.380 50.360 ;
        RECT 117.500 50.040 117.820 50.360 ;
        RECT 4.180 48.640 4.500 48.960 ;
        RECT 4.620 48.640 4.940 48.960 ;
        RECT 5.060 48.640 5.380 48.960 ;
        RECT 5.500 48.640 5.820 48.960 ;
        RECT 32.180 24.890 32.500 25.210 ;
        RECT 32.620 24.890 32.940 25.210 ;
        RECT 33.060 24.890 33.380 25.210 ;
        RECT 33.500 24.890 33.820 25.210 ;
        RECT 60.180 24.890 60.500 25.210 ;
        RECT 60.620 24.890 60.940 25.210 ;
        RECT 61.060 24.890 61.380 25.210 ;
        RECT 61.500 24.890 61.820 25.210 ;
      LAYER met3 ;
        RECT 4.000 87.000 118.000 89.000 ;
        RECT 32.000 56.610 34.000 57.090 ;
        RECT 60.000 56.610 62.000 57.090 ;
        RECT 88.000 56.610 90.000 57.090 ;
        RECT 116.000 49.960 118.000 50.440 ;
        RECT 4.000 48.560 6.000 49.040 ;
        RECT 32.000 24.810 34.000 25.290 ;
        RECT 60.000 24.810 62.000 25.290 ;
        RECT 4.000 -8.000 118.000 -6.000 ;
      LAYER via3 ;
        RECT 4.200 88.400 4.600 88.800 ;
        RECT 4.800 88.400 5.200 88.800 ;
        RECT 5.400 88.400 5.800 88.800 ;
        RECT 32.200 88.400 32.600 88.800 ;
        RECT 32.800 88.400 33.200 88.800 ;
        RECT 33.400 88.400 33.800 88.800 ;
        RECT 60.200 88.400 60.600 88.800 ;
        RECT 60.800 88.400 61.200 88.800 ;
        RECT 61.400 88.400 61.800 88.800 ;
        RECT 88.200 88.400 88.600 88.800 ;
        RECT 88.800 88.400 89.200 88.800 ;
        RECT 89.400 88.400 89.800 88.800 ;
        RECT 116.200 88.400 116.600 88.800 ;
        RECT 116.800 88.400 117.200 88.800 ;
        RECT 117.400 88.400 117.800 88.800 ;
        RECT 4.200 87.800 4.600 88.200 ;
        RECT 4.800 87.800 5.200 88.200 ;
        RECT 5.400 87.800 5.800 88.200 ;
        RECT 32.200 87.800 32.600 88.200 ;
        RECT 32.800 87.800 33.200 88.200 ;
        RECT 33.400 87.800 33.800 88.200 ;
        RECT 60.200 87.800 60.600 88.200 ;
        RECT 60.800 87.800 61.200 88.200 ;
        RECT 61.400 87.800 61.800 88.200 ;
        RECT 88.200 87.800 88.600 88.200 ;
        RECT 88.800 87.800 89.200 88.200 ;
        RECT 89.400 87.800 89.800 88.200 ;
        RECT 116.200 87.800 116.600 88.200 ;
        RECT 116.800 87.800 117.200 88.200 ;
        RECT 117.400 87.800 117.800 88.200 ;
        RECT 4.200 87.200 4.600 87.600 ;
        RECT 4.800 87.200 5.200 87.600 ;
        RECT 5.400 87.200 5.800 87.600 ;
        RECT 32.200 87.200 32.600 87.600 ;
        RECT 32.800 87.200 33.200 87.600 ;
        RECT 33.400 87.200 33.800 87.600 ;
        RECT 60.200 87.200 60.600 87.600 ;
        RECT 60.800 87.200 61.200 87.600 ;
        RECT 61.400 87.200 61.800 87.600 ;
        RECT 88.200 87.200 88.600 87.600 ;
        RECT 88.800 87.200 89.200 87.600 ;
        RECT 89.400 87.200 89.800 87.600 ;
        RECT 116.200 87.200 116.600 87.600 ;
        RECT 116.800 87.200 117.200 87.600 ;
        RECT 117.400 87.200 117.800 87.600 ;
        RECT 32.160 56.670 32.520 57.035 ;
        RECT 32.600 56.670 32.960 57.035 ;
        RECT 33.040 56.670 33.400 57.035 ;
        RECT 33.480 56.670 33.840 57.035 ;
        RECT 60.160 56.670 60.520 57.035 ;
        RECT 60.600 56.670 60.960 57.035 ;
        RECT 61.040 56.670 61.400 57.035 ;
        RECT 61.480 56.670 61.840 57.035 ;
        RECT 88.160 56.670 88.520 57.035 ;
        RECT 88.600 56.670 88.960 57.035 ;
        RECT 89.040 56.670 89.400 57.035 ;
        RECT 89.480 56.670 89.840 57.035 ;
        RECT 116.160 50.020 116.520 50.385 ;
        RECT 116.600 50.020 116.960 50.385 ;
        RECT 117.040 50.020 117.400 50.385 ;
        RECT 117.480 50.020 117.840 50.385 ;
        RECT 4.160 48.620 4.520 48.985 ;
        RECT 4.600 48.620 4.960 48.985 ;
        RECT 5.040 48.620 5.400 48.985 ;
        RECT 5.480 48.620 5.840 48.985 ;
        RECT 32.160 24.870 32.520 25.235 ;
        RECT 32.600 24.870 32.960 25.235 ;
        RECT 33.040 24.870 33.400 25.235 ;
        RECT 33.480 24.870 33.840 25.235 ;
        RECT 60.160 24.870 60.520 25.235 ;
        RECT 60.600 24.870 60.960 25.235 ;
        RECT 61.040 24.870 61.400 25.235 ;
        RECT 61.480 24.870 61.840 25.235 ;
        RECT 4.200 -6.600 4.600 -6.200 ;
        RECT 4.800 -6.600 5.200 -6.200 ;
        RECT 5.400 -6.600 5.800 -6.200 ;
        RECT 32.200 -6.600 32.600 -6.200 ;
        RECT 32.800 -6.600 33.200 -6.200 ;
        RECT 33.400 -6.600 33.800 -6.200 ;
        RECT 60.200 -6.600 60.600 -6.200 ;
        RECT 60.800 -6.600 61.200 -6.200 ;
        RECT 61.400 -6.600 61.800 -6.200 ;
        RECT 88.200 -6.600 88.600 -6.200 ;
        RECT 88.800 -6.600 89.200 -6.200 ;
        RECT 89.400 -6.600 89.800 -6.200 ;
        RECT 116.200 -6.600 116.600 -6.200 ;
        RECT 116.800 -6.600 117.200 -6.200 ;
        RECT 117.400 -6.600 117.800 -6.200 ;
        RECT 4.200 -7.200 4.600 -6.800 ;
        RECT 4.800 -7.200 5.200 -6.800 ;
        RECT 5.400 -7.200 5.800 -6.800 ;
        RECT 32.200 -7.200 32.600 -6.800 ;
        RECT 32.800 -7.200 33.200 -6.800 ;
        RECT 33.400 -7.200 33.800 -6.800 ;
        RECT 60.200 -7.200 60.600 -6.800 ;
        RECT 60.800 -7.200 61.200 -6.800 ;
        RECT 61.400 -7.200 61.800 -6.800 ;
        RECT 88.200 -7.200 88.600 -6.800 ;
        RECT 88.800 -7.200 89.200 -6.800 ;
        RECT 89.400 -7.200 89.800 -6.800 ;
        RECT 116.200 -7.200 116.600 -6.800 ;
        RECT 116.800 -7.200 117.200 -6.800 ;
        RECT 117.400 -7.200 117.800 -6.800 ;
        RECT 4.200 -7.800 4.600 -7.400 ;
        RECT 4.800 -7.800 5.200 -7.400 ;
        RECT 5.400 -7.800 5.800 -7.400 ;
        RECT 32.200 -7.800 32.600 -7.400 ;
        RECT 32.800 -7.800 33.200 -7.400 ;
        RECT 33.400 -7.800 33.800 -7.400 ;
        RECT 60.200 -7.800 60.600 -7.400 ;
        RECT 60.800 -7.800 61.200 -7.400 ;
        RECT 61.400 -7.800 61.800 -7.400 ;
        RECT 88.200 -7.800 88.600 -7.400 ;
        RECT 88.800 -7.800 89.200 -7.400 ;
        RECT 89.400 -7.800 89.800 -7.400 ;
        RECT 116.200 -7.800 116.600 -7.400 ;
        RECT 116.800 -7.800 117.200 -7.400 ;
        RECT 117.400 -7.800 117.800 -7.400 ;
      LAYER met4 ;
        RECT 4.000 -8.000 6.000 89.000 ;
        RECT 32.000 -8.000 34.000 89.000 ;
        RECT 60.000 -8.000 62.000 89.000 ;
        RECT 88.000 -8.000 90.000 89.000 ;
        RECT 116.000 -8.000 118.000 89.000 ;
    END
  END vssd2
  OBS
      LAYER pwell ;
        RECT 7.180 49.585 8.985 49.815 ;
        RECT 6.695 48.905 8.985 49.585 ;
        RECT 6.840 48.715 7.010 48.905 ;
        RECT 10.830 48.715 11.000 48.885 ;
        RECT 15.980 41.470 105.050 48.570 ;
        RECT 108.000 46.000 111.000 51.000 ;
        RECT 108.000 45.000 116.000 46.000 ;
        RECT 110.000 43.000 116.000 45.000 ;
        RECT 7.500 33.270 114.280 40.370 ;
      LAYER li1 ;
        RECT 6.775 50.865 7.035 51.265 ;
        RECT 6.775 50.695 8.140 50.865 ;
        RECT 7.405 49.625 8.140 50.695 ;
        RECT 8.665 50.750 8.905 50.755 ;
        RECT 9.180 50.750 10.505 50.960 ;
        RECT 8.665 50.740 10.505 50.750 ;
        RECT 8.665 50.530 9.400 50.740 ;
        RECT 10.285 50.535 10.505 50.740 ;
        RECT 10.770 50.535 11.290 50.540 ;
        RECT 8.665 49.775 8.905 50.530 ;
        RECT 10.285 50.315 11.290 50.535 ;
        RECT 6.775 49.455 8.140 49.625 ;
        RECT 6.775 49.055 7.035 49.455 ;
        RECT 10.770 49.055 11.290 50.315 ;
        RECT 11.460 49.715 11.980 51.265 ;
        RECT 23.400 48.950 23.780 49.000 ;
        RECT 22.450 48.590 23.780 48.950 ;
        RECT 23.400 48.540 23.780 48.590 ;
        RECT 16.670 42.090 16.960 47.540 ;
        RECT 21.050 42.090 21.340 47.540 ;
        RECT 22.190 42.090 22.480 47.540 ;
        RECT 24.375 42.500 24.675 55.090 ;
        RECT 25.270 48.950 25.650 49.000 ;
        RECT 25.270 48.590 26.600 48.950 ;
        RECT 25.270 48.540 25.650 48.590 ;
        RECT 26.570 42.090 26.860 47.540 ;
        RECT 27.710 42.090 28.000 47.540 ;
        RECT 29.900 42.500 30.200 55.090 ;
        RECT 32.250 48.950 32.630 49.000 ;
        RECT 41.110 48.950 41.490 49.000 ;
        RECT 31.300 48.590 32.630 48.950 ;
        RECT 40.160 48.590 41.490 48.950 ;
        RECT 32.250 48.540 32.630 48.590 ;
        RECT 41.110 48.540 41.490 48.590 ;
        RECT 31.040 42.090 31.330 47.540 ;
        RECT 34.380 42.090 34.670 47.540 ;
        RECT 38.760 42.090 39.050 47.540 ;
        RECT 39.900 42.090 40.190 47.540 ;
        RECT 42.085 42.500 42.385 55.090 ;
        RECT 42.980 48.950 43.360 49.000 ;
        RECT 42.980 48.590 44.310 48.950 ;
        RECT 42.980 48.540 43.360 48.590 ;
        RECT 44.280 42.090 44.570 47.540 ;
        RECT 45.420 42.090 45.710 47.540 ;
        RECT 47.610 42.500 47.910 55.090 ;
        RECT 49.960 48.950 50.340 49.000 ;
        RECT 58.820 48.950 59.200 49.000 ;
        RECT 49.010 48.590 50.340 48.950 ;
        RECT 57.870 48.590 59.200 48.950 ;
        RECT 49.960 48.540 50.340 48.590 ;
        RECT 58.820 48.540 59.200 48.590 ;
        RECT 48.750 42.090 49.040 47.540 ;
        RECT 52.090 42.090 52.380 47.540 ;
        RECT 56.470 42.090 56.760 47.540 ;
        RECT 57.610 42.090 57.900 47.540 ;
        RECT 59.795 42.500 60.095 55.090 ;
        RECT 60.690 48.950 61.070 49.000 ;
        RECT 60.690 48.590 62.020 48.950 ;
        RECT 60.690 48.540 61.070 48.590 ;
        RECT 61.990 42.090 62.280 47.540 ;
        RECT 63.130 42.090 63.420 47.540 ;
        RECT 65.320 42.500 65.620 55.090 ;
        RECT 67.670 48.950 68.050 49.000 ;
        RECT 76.530 48.950 76.910 49.000 ;
        RECT 66.720 48.590 68.050 48.950 ;
        RECT 75.580 48.590 76.910 48.950 ;
        RECT 67.670 48.540 68.050 48.590 ;
        RECT 76.530 48.540 76.910 48.590 ;
        RECT 66.460 42.090 66.750 47.540 ;
        RECT 69.800 42.090 70.090 47.540 ;
        RECT 74.180 42.090 74.470 47.540 ;
        RECT 75.320 42.090 75.610 47.540 ;
        RECT 77.505 42.500 77.805 55.090 ;
        RECT 78.400 48.950 78.780 49.000 ;
        RECT 78.400 48.590 79.730 48.950 ;
        RECT 78.400 48.540 78.780 48.590 ;
        RECT 79.700 42.090 79.990 47.540 ;
        RECT 80.840 42.090 81.130 47.540 ;
        RECT 83.030 42.500 83.330 55.090 ;
        RECT 85.380 48.950 85.760 49.000 ;
        RECT 94.240 48.950 94.620 49.000 ;
        RECT 84.430 48.590 85.760 48.950 ;
        RECT 93.290 48.590 94.620 48.950 ;
        RECT 85.380 48.540 85.760 48.590 ;
        RECT 94.240 48.540 94.620 48.590 ;
        RECT 84.170 42.090 84.460 47.540 ;
        RECT 87.510 42.090 87.800 47.540 ;
        RECT 91.890 42.090 92.180 47.540 ;
        RECT 93.030 42.090 93.320 47.540 ;
        RECT 95.215 42.500 95.515 55.090 ;
        RECT 96.110 48.950 96.490 49.000 ;
        RECT 96.110 48.590 97.440 48.950 ;
        RECT 96.110 48.540 96.490 48.590 ;
        RECT 97.410 42.090 97.700 47.540 ;
        RECT 98.550 42.090 98.840 47.540 ;
        RECT 100.740 42.500 101.040 55.090 ;
        RECT 103.090 48.950 103.470 49.000 ;
        RECT 102.140 48.590 103.470 48.950 ;
        RECT 103.090 48.540 103.470 48.590 ;
        RECT 101.880 42.090 102.170 47.540 ;
        RECT 108.500 45.500 110.500 45.865 ;
        RECT 109.500 44.500 110.865 45.500 ;
        RECT 110.500 43.500 110.865 44.500 ;
        RECT 16.160 41.730 18.050 42.090 ;
        RECT 19.840 41.730 23.690 42.090 ;
        RECT 25.350 41.730 29.200 42.090 ;
        RECT 31.040 41.730 32.440 42.090 ;
        RECT 33.870 41.730 35.760 42.090 ;
        RECT 37.550 41.730 41.400 42.090 ;
        RECT 43.060 41.730 46.910 42.090 ;
        RECT 48.750 41.730 50.150 42.090 ;
        RECT 51.580 41.730 53.470 42.090 ;
        RECT 55.260 41.730 59.110 42.090 ;
        RECT 60.770 41.730 64.620 42.090 ;
        RECT 66.460 41.730 67.860 42.090 ;
        RECT 69.290 41.730 71.180 42.090 ;
        RECT 72.970 41.730 76.820 42.090 ;
        RECT 78.480 41.730 82.330 42.090 ;
        RECT 84.170 41.730 85.570 42.090 ;
        RECT 87.000 41.730 88.890 42.090 ;
        RECT 90.680 41.730 94.530 42.090 ;
        RECT 96.190 41.730 100.040 42.090 ;
        RECT 101.880 41.730 103.280 42.090 ;
        RECT 9.270 39.750 10.670 40.110 ;
        RECT 12.510 39.750 16.360 40.110 ;
        RECT 18.020 39.750 21.870 40.110 ;
        RECT 23.660 39.750 25.550 40.110 ;
        RECT 26.980 39.750 28.380 40.110 ;
        RECT 30.220 39.750 34.070 40.110 ;
        RECT 35.730 39.750 39.580 40.110 ;
        RECT 41.370 39.750 43.260 40.110 ;
        RECT 44.690 39.750 46.090 40.110 ;
        RECT 47.930 39.750 51.780 40.110 ;
        RECT 53.440 39.750 57.290 40.110 ;
        RECT 59.080 39.750 60.970 40.110 ;
        RECT 62.400 39.750 63.800 40.110 ;
        RECT 65.640 39.750 69.490 40.110 ;
        RECT 71.150 39.750 75.000 40.110 ;
        RECT 76.790 39.750 78.680 40.110 ;
        RECT 80.110 39.750 81.510 40.110 ;
        RECT 83.350 39.750 87.200 40.110 ;
        RECT 88.860 39.750 92.710 40.110 ;
        RECT 94.500 39.750 96.390 40.110 ;
        RECT 97.820 39.750 99.220 40.110 ;
        RECT 101.060 39.750 104.910 40.110 ;
        RECT 106.570 39.750 110.420 40.110 ;
        RECT 112.210 39.750 114.100 40.110 ;
        RECT 10.380 34.300 10.670 39.750 ;
        RECT 9.080 33.250 9.460 33.300 ;
        RECT 9.080 32.890 10.410 33.250 ;
        RECT 9.080 32.840 9.460 32.890 ;
        RECT 11.510 26.750 11.810 39.340 ;
        RECT 13.710 34.300 14.000 39.750 ;
        RECT 14.850 34.300 15.140 39.750 ;
        RECT 16.060 33.250 16.440 33.300 ;
        RECT 15.110 32.890 16.440 33.250 ;
        RECT 16.060 32.840 16.440 32.890 ;
        RECT 17.035 26.750 17.335 39.340 ;
        RECT 19.230 34.300 19.520 39.750 ;
        RECT 20.370 34.300 20.660 39.750 ;
        RECT 24.750 34.300 25.040 39.750 ;
        RECT 28.090 34.300 28.380 39.750 ;
        RECT 17.930 33.250 18.310 33.300 ;
        RECT 26.790 33.250 27.170 33.300 ;
        RECT 17.930 32.890 19.260 33.250 ;
        RECT 26.790 32.890 28.120 33.250 ;
        RECT 17.930 32.840 18.310 32.890 ;
        RECT 26.790 32.840 27.170 32.890 ;
        RECT 29.220 26.750 29.520 39.340 ;
        RECT 31.420 34.300 31.710 39.750 ;
        RECT 32.560 34.300 32.850 39.750 ;
        RECT 33.770 33.250 34.150 33.300 ;
        RECT 32.820 32.890 34.150 33.250 ;
        RECT 33.770 32.840 34.150 32.890 ;
        RECT 34.745 26.750 35.045 39.340 ;
        RECT 36.940 34.300 37.230 39.750 ;
        RECT 38.080 34.300 38.370 39.750 ;
        RECT 42.460 34.300 42.750 39.750 ;
        RECT 45.800 34.300 46.090 39.750 ;
        RECT 35.640 33.250 36.020 33.300 ;
        RECT 44.500 33.250 44.880 33.300 ;
        RECT 35.640 32.890 36.970 33.250 ;
        RECT 44.500 32.890 45.830 33.250 ;
        RECT 35.640 32.840 36.020 32.890 ;
        RECT 44.500 32.840 44.880 32.890 ;
        RECT 46.930 26.750 47.230 39.340 ;
        RECT 49.130 34.300 49.420 39.750 ;
        RECT 50.270 34.300 50.560 39.750 ;
        RECT 51.480 33.250 51.860 33.300 ;
        RECT 50.530 32.890 51.860 33.250 ;
        RECT 51.480 32.840 51.860 32.890 ;
        RECT 52.455 26.750 52.755 39.340 ;
        RECT 54.650 34.300 54.940 39.750 ;
        RECT 55.790 34.300 56.080 39.750 ;
        RECT 60.170 34.300 60.460 39.750 ;
        RECT 63.510 34.300 63.800 39.750 ;
        RECT 53.350 33.250 53.730 33.300 ;
        RECT 62.210 33.250 62.590 33.300 ;
        RECT 53.350 32.890 54.680 33.250 ;
        RECT 62.210 32.890 63.540 33.250 ;
        RECT 53.350 32.840 53.730 32.890 ;
        RECT 62.210 32.840 62.590 32.890 ;
        RECT 64.640 26.750 64.940 39.340 ;
        RECT 66.840 34.300 67.130 39.750 ;
        RECT 67.980 34.300 68.270 39.750 ;
        RECT 69.190 33.250 69.570 33.300 ;
        RECT 68.240 32.890 69.570 33.250 ;
        RECT 69.190 32.840 69.570 32.890 ;
        RECT 70.165 26.750 70.465 39.340 ;
        RECT 72.360 34.300 72.650 39.750 ;
        RECT 73.500 34.300 73.790 39.750 ;
        RECT 77.880 34.300 78.170 39.750 ;
        RECT 81.220 34.300 81.510 39.750 ;
        RECT 71.060 33.250 71.440 33.300 ;
        RECT 79.920 33.250 80.300 33.300 ;
        RECT 71.060 32.890 72.390 33.250 ;
        RECT 79.920 32.890 81.250 33.250 ;
        RECT 71.060 32.840 71.440 32.890 ;
        RECT 79.920 32.840 80.300 32.890 ;
        RECT 82.350 26.750 82.650 39.340 ;
        RECT 84.550 34.300 84.840 39.750 ;
        RECT 85.690 34.300 85.980 39.750 ;
        RECT 86.900 33.250 87.280 33.300 ;
        RECT 85.950 32.890 87.280 33.250 ;
        RECT 86.900 32.840 87.280 32.890 ;
        RECT 87.875 26.750 88.175 39.340 ;
        RECT 90.070 34.300 90.360 39.750 ;
        RECT 91.210 34.300 91.500 39.750 ;
        RECT 95.590 34.300 95.880 39.750 ;
        RECT 98.930 34.300 99.220 39.750 ;
        RECT 88.770 33.250 89.150 33.300 ;
        RECT 97.630 33.250 98.010 33.300 ;
        RECT 88.770 32.890 90.100 33.250 ;
        RECT 97.630 32.890 98.960 33.250 ;
        RECT 88.770 32.840 89.150 32.890 ;
        RECT 97.630 32.840 98.010 32.890 ;
        RECT 100.060 26.750 100.360 39.340 ;
        RECT 102.260 34.300 102.550 39.750 ;
        RECT 103.400 34.300 103.690 39.750 ;
        RECT 104.610 33.250 104.990 33.300 ;
        RECT 103.660 32.890 104.990 33.250 ;
        RECT 104.610 32.840 104.990 32.890 ;
        RECT 105.585 26.750 105.885 39.340 ;
        RECT 107.780 34.300 108.070 39.750 ;
        RECT 108.920 34.300 109.210 39.750 ;
        RECT 113.300 34.300 113.590 39.750 ;
        RECT 106.480 33.250 106.860 33.300 ;
        RECT 106.480 32.890 107.810 33.250 ;
        RECT 106.480 32.840 106.860 32.890 ;
      LAYER mcon ;
        RECT 22.450 48.620 22.750 48.920 ;
        RECT 22.940 48.620 23.240 48.920 ;
        RECT 23.430 48.620 23.730 48.920 ;
        RECT 25.320 48.620 25.620 48.920 ;
        RECT 25.810 48.620 26.110 48.920 ;
        RECT 26.300 48.620 26.600 48.920 ;
        RECT 24.375 47.260 24.675 47.560 ;
        RECT 31.300 48.620 31.600 48.920 ;
        RECT 31.790 48.620 32.090 48.920 ;
        RECT 32.280 48.620 32.580 48.920 ;
        RECT 40.160 48.620 40.460 48.920 ;
        RECT 40.650 48.620 40.950 48.920 ;
        RECT 41.140 48.620 41.440 48.920 ;
        RECT 29.900 47.260 30.200 47.560 ;
        RECT 43.030 48.620 43.330 48.920 ;
        RECT 43.520 48.620 43.820 48.920 ;
        RECT 44.010 48.620 44.310 48.920 ;
        RECT 42.085 47.260 42.385 47.560 ;
        RECT 49.010 48.620 49.310 48.920 ;
        RECT 49.500 48.620 49.800 48.920 ;
        RECT 49.990 48.620 50.290 48.920 ;
        RECT 57.870 48.620 58.170 48.920 ;
        RECT 58.360 48.620 58.660 48.920 ;
        RECT 58.850 48.620 59.150 48.920 ;
        RECT 47.610 47.260 47.910 47.560 ;
        RECT 60.740 48.620 61.040 48.920 ;
        RECT 61.230 48.620 61.530 48.920 ;
        RECT 61.720 48.620 62.020 48.920 ;
        RECT 59.795 47.260 60.095 47.560 ;
        RECT 66.720 48.620 67.020 48.920 ;
        RECT 67.210 48.620 67.510 48.920 ;
        RECT 67.700 48.620 68.000 48.920 ;
        RECT 75.580 48.620 75.880 48.920 ;
        RECT 76.070 48.620 76.370 48.920 ;
        RECT 76.560 48.620 76.860 48.920 ;
        RECT 65.320 47.260 65.620 47.560 ;
        RECT 78.450 48.620 78.750 48.920 ;
        RECT 78.940 48.620 79.240 48.920 ;
        RECT 79.430 48.620 79.730 48.920 ;
        RECT 77.505 47.260 77.805 47.560 ;
        RECT 84.430 48.620 84.730 48.920 ;
        RECT 84.920 48.620 85.220 48.920 ;
        RECT 85.410 48.620 85.710 48.920 ;
        RECT 93.290 48.620 93.590 48.920 ;
        RECT 93.780 48.620 94.080 48.920 ;
        RECT 94.270 48.620 94.570 48.920 ;
        RECT 83.030 47.260 83.330 47.560 ;
        RECT 96.160 48.620 96.460 48.920 ;
        RECT 96.650 48.620 96.950 48.920 ;
        RECT 97.140 48.620 97.440 48.920 ;
        RECT 95.215 47.260 95.515 47.560 ;
        RECT 102.140 48.620 102.440 48.920 ;
        RECT 102.630 48.620 102.930 48.920 ;
        RECT 103.120 48.620 103.420 48.920 ;
        RECT 100.740 47.260 101.040 47.560 ;
        RECT 109.590 45.120 109.890 45.420 ;
        RECT 110.110 45.120 110.410 45.420 ;
        RECT 109.590 44.600 109.890 44.900 ;
        RECT 110.110 44.600 110.410 44.900 ;
        RECT 16.220 41.760 16.520 42.060 ;
        RECT 16.710 41.760 17.010 42.060 ;
        RECT 17.200 41.760 17.500 42.060 ;
        RECT 17.690 41.760 17.990 42.060 ;
        RECT 19.900 41.760 20.200 42.060 ;
        RECT 20.390 41.760 20.690 42.060 ;
        RECT 20.880 41.760 21.180 42.060 ;
        RECT 21.370 41.760 21.670 42.060 ;
        RECT 21.860 41.760 22.160 42.060 ;
        RECT 22.350 41.760 22.650 42.060 ;
        RECT 22.840 41.760 23.140 42.060 ;
        RECT 23.330 41.760 23.630 42.060 ;
        RECT 25.410 41.760 25.710 42.060 ;
        RECT 25.900 41.760 26.200 42.060 ;
        RECT 26.390 41.760 26.690 42.060 ;
        RECT 26.880 41.760 27.180 42.060 ;
        RECT 27.370 41.760 27.670 42.060 ;
        RECT 27.860 41.760 28.160 42.060 ;
        RECT 28.350 41.760 28.650 42.060 ;
        RECT 28.840 41.760 29.140 42.060 ;
        RECT 31.100 41.760 31.400 42.060 ;
        RECT 31.590 41.760 31.890 42.060 ;
        RECT 32.080 41.760 32.380 42.060 ;
        RECT 33.930 41.760 34.230 42.060 ;
        RECT 34.420 41.760 34.720 42.060 ;
        RECT 34.910 41.760 35.210 42.060 ;
        RECT 35.400 41.760 35.700 42.060 ;
        RECT 37.610 41.760 37.910 42.060 ;
        RECT 38.100 41.760 38.400 42.060 ;
        RECT 38.590 41.760 38.890 42.060 ;
        RECT 39.080 41.760 39.380 42.060 ;
        RECT 39.570 41.760 39.870 42.060 ;
        RECT 40.060 41.760 40.360 42.060 ;
        RECT 40.550 41.760 40.850 42.060 ;
        RECT 41.040 41.760 41.340 42.060 ;
        RECT 43.120 41.760 43.420 42.060 ;
        RECT 43.610 41.760 43.910 42.060 ;
        RECT 44.100 41.760 44.400 42.060 ;
        RECT 44.590 41.760 44.890 42.060 ;
        RECT 45.080 41.760 45.380 42.060 ;
        RECT 45.570 41.760 45.870 42.060 ;
        RECT 46.060 41.760 46.360 42.060 ;
        RECT 46.550 41.760 46.850 42.060 ;
        RECT 48.810 41.760 49.110 42.060 ;
        RECT 49.300 41.760 49.600 42.060 ;
        RECT 49.790 41.760 50.090 42.060 ;
        RECT 51.640 41.760 51.940 42.060 ;
        RECT 52.130 41.760 52.430 42.060 ;
        RECT 52.620 41.760 52.920 42.060 ;
        RECT 53.110 41.760 53.410 42.060 ;
        RECT 55.320 41.760 55.620 42.060 ;
        RECT 55.810 41.760 56.110 42.060 ;
        RECT 56.300 41.760 56.600 42.060 ;
        RECT 56.790 41.760 57.090 42.060 ;
        RECT 57.280 41.760 57.580 42.060 ;
        RECT 57.770 41.760 58.070 42.060 ;
        RECT 58.260 41.760 58.560 42.060 ;
        RECT 58.750 41.760 59.050 42.060 ;
        RECT 60.830 41.760 61.130 42.060 ;
        RECT 61.320 41.760 61.620 42.060 ;
        RECT 61.810 41.760 62.110 42.060 ;
        RECT 62.300 41.760 62.600 42.060 ;
        RECT 62.790 41.760 63.090 42.060 ;
        RECT 63.280 41.760 63.580 42.060 ;
        RECT 63.770 41.760 64.070 42.060 ;
        RECT 64.260 41.760 64.560 42.060 ;
        RECT 66.520 41.760 66.820 42.060 ;
        RECT 67.010 41.760 67.310 42.060 ;
        RECT 67.500 41.760 67.800 42.060 ;
        RECT 69.350 41.760 69.650 42.060 ;
        RECT 69.840 41.760 70.140 42.060 ;
        RECT 70.330 41.760 70.630 42.060 ;
        RECT 70.820 41.760 71.120 42.060 ;
        RECT 73.030 41.760 73.330 42.060 ;
        RECT 73.520 41.760 73.820 42.060 ;
        RECT 74.010 41.760 74.310 42.060 ;
        RECT 74.500 41.760 74.800 42.060 ;
        RECT 74.990 41.760 75.290 42.060 ;
        RECT 75.480 41.760 75.780 42.060 ;
        RECT 75.970 41.760 76.270 42.060 ;
        RECT 76.460 41.760 76.760 42.060 ;
        RECT 78.540 41.760 78.840 42.060 ;
        RECT 79.030 41.760 79.330 42.060 ;
        RECT 79.520 41.760 79.820 42.060 ;
        RECT 80.010 41.760 80.310 42.060 ;
        RECT 80.500 41.760 80.800 42.060 ;
        RECT 80.990 41.760 81.290 42.060 ;
        RECT 81.480 41.760 81.780 42.060 ;
        RECT 81.970 41.760 82.270 42.060 ;
        RECT 84.230 41.760 84.530 42.060 ;
        RECT 84.720 41.760 85.020 42.060 ;
        RECT 85.210 41.760 85.510 42.060 ;
        RECT 87.060 41.760 87.360 42.060 ;
        RECT 87.550 41.760 87.850 42.060 ;
        RECT 88.040 41.760 88.340 42.060 ;
        RECT 88.530 41.760 88.830 42.060 ;
        RECT 90.740 41.760 91.040 42.060 ;
        RECT 91.230 41.760 91.530 42.060 ;
        RECT 91.720 41.760 92.020 42.060 ;
        RECT 92.210 41.760 92.510 42.060 ;
        RECT 92.700 41.760 93.000 42.060 ;
        RECT 93.190 41.760 93.490 42.060 ;
        RECT 93.680 41.760 93.980 42.060 ;
        RECT 94.170 41.760 94.470 42.060 ;
        RECT 96.250 41.760 96.550 42.060 ;
        RECT 96.740 41.760 97.040 42.060 ;
        RECT 97.230 41.760 97.530 42.060 ;
        RECT 97.720 41.760 98.020 42.060 ;
        RECT 98.210 41.760 98.510 42.060 ;
        RECT 98.700 41.760 99.000 42.060 ;
        RECT 99.190 41.760 99.490 42.060 ;
        RECT 99.680 41.760 99.980 42.060 ;
        RECT 101.940 41.760 102.240 42.060 ;
        RECT 102.430 41.760 102.730 42.060 ;
        RECT 102.920 41.760 103.220 42.060 ;
        RECT 9.330 39.780 9.630 40.080 ;
        RECT 9.820 39.780 10.120 40.080 ;
        RECT 10.310 39.780 10.610 40.080 ;
        RECT 12.570 39.780 12.870 40.080 ;
        RECT 13.060 39.780 13.360 40.080 ;
        RECT 13.550 39.780 13.850 40.080 ;
        RECT 14.040 39.780 14.340 40.080 ;
        RECT 14.530 39.780 14.830 40.080 ;
        RECT 15.020 39.780 15.320 40.080 ;
        RECT 15.510 39.780 15.810 40.080 ;
        RECT 16.000 39.780 16.300 40.080 ;
        RECT 18.080 39.780 18.380 40.080 ;
        RECT 18.570 39.780 18.870 40.080 ;
        RECT 19.060 39.780 19.360 40.080 ;
        RECT 19.550 39.780 19.850 40.080 ;
        RECT 20.040 39.780 20.340 40.080 ;
        RECT 20.530 39.780 20.830 40.080 ;
        RECT 21.020 39.780 21.320 40.080 ;
        RECT 21.510 39.780 21.810 40.080 ;
        RECT 23.720 39.780 24.020 40.080 ;
        RECT 24.210 39.780 24.510 40.080 ;
        RECT 24.700 39.780 25.000 40.080 ;
        RECT 25.190 39.780 25.490 40.080 ;
        RECT 27.040 39.780 27.340 40.080 ;
        RECT 27.530 39.780 27.830 40.080 ;
        RECT 28.020 39.780 28.320 40.080 ;
        RECT 30.280 39.780 30.580 40.080 ;
        RECT 30.770 39.780 31.070 40.080 ;
        RECT 31.260 39.780 31.560 40.080 ;
        RECT 31.750 39.780 32.050 40.080 ;
        RECT 32.240 39.780 32.540 40.080 ;
        RECT 32.730 39.780 33.030 40.080 ;
        RECT 33.220 39.780 33.520 40.080 ;
        RECT 33.710 39.780 34.010 40.080 ;
        RECT 35.790 39.780 36.090 40.080 ;
        RECT 36.280 39.780 36.580 40.080 ;
        RECT 36.770 39.780 37.070 40.080 ;
        RECT 37.260 39.780 37.560 40.080 ;
        RECT 37.750 39.780 38.050 40.080 ;
        RECT 38.240 39.780 38.540 40.080 ;
        RECT 38.730 39.780 39.030 40.080 ;
        RECT 39.220 39.780 39.520 40.080 ;
        RECT 41.430 39.780 41.730 40.080 ;
        RECT 41.920 39.780 42.220 40.080 ;
        RECT 42.410 39.780 42.710 40.080 ;
        RECT 42.900 39.780 43.200 40.080 ;
        RECT 44.750 39.780 45.050 40.080 ;
        RECT 45.240 39.780 45.540 40.080 ;
        RECT 45.730 39.780 46.030 40.080 ;
        RECT 47.990 39.780 48.290 40.080 ;
        RECT 48.480 39.780 48.780 40.080 ;
        RECT 48.970 39.780 49.270 40.080 ;
        RECT 49.460 39.780 49.760 40.080 ;
        RECT 49.950 39.780 50.250 40.080 ;
        RECT 50.440 39.780 50.740 40.080 ;
        RECT 50.930 39.780 51.230 40.080 ;
        RECT 51.420 39.780 51.720 40.080 ;
        RECT 53.500 39.780 53.800 40.080 ;
        RECT 53.990 39.780 54.290 40.080 ;
        RECT 54.480 39.780 54.780 40.080 ;
        RECT 54.970 39.780 55.270 40.080 ;
        RECT 55.460 39.780 55.760 40.080 ;
        RECT 55.950 39.780 56.250 40.080 ;
        RECT 56.440 39.780 56.740 40.080 ;
        RECT 56.930 39.780 57.230 40.080 ;
        RECT 59.140 39.780 59.440 40.080 ;
        RECT 59.630 39.780 59.930 40.080 ;
        RECT 60.120 39.780 60.420 40.080 ;
        RECT 60.610 39.780 60.910 40.080 ;
        RECT 62.460 39.780 62.760 40.080 ;
        RECT 62.950 39.780 63.250 40.080 ;
        RECT 63.440 39.780 63.740 40.080 ;
        RECT 65.700 39.780 66.000 40.080 ;
        RECT 66.190 39.780 66.490 40.080 ;
        RECT 66.680 39.780 66.980 40.080 ;
        RECT 67.170 39.780 67.470 40.080 ;
        RECT 67.660 39.780 67.960 40.080 ;
        RECT 68.150 39.780 68.450 40.080 ;
        RECT 68.640 39.780 68.940 40.080 ;
        RECT 69.130 39.780 69.430 40.080 ;
        RECT 71.210 39.780 71.510 40.080 ;
        RECT 71.700 39.780 72.000 40.080 ;
        RECT 72.190 39.780 72.490 40.080 ;
        RECT 72.680 39.780 72.980 40.080 ;
        RECT 73.170 39.780 73.470 40.080 ;
        RECT 73.660 39.780 73.960 40.080 ;
        RECT 74.150 39.780 74.450 40.080 ;
        RECT 74.640 39.780 74.940 40.080 ;
        RECT 76.850 39.780 77.150 40.080 ;
        RECT 77.340 39.780 77.640 40.080 ;
        RECT 77.830 39.780 78.130 40.080 ;
        RECT 78.320 39.780 78.620 40.080 ;
        RECT 80.170 39.780 80.470 40.080 ;
        RECT 80.660 39.780 80.960 40.080 ;
        RECT 81.150 39.780 81.450 40.080 ;
        RECT 83.410 39.780 83.710 40.080 ;
        RECT 83.900 39.780 84.200 40.080 ;
        RECT 84.390 39.780 84.690 40.080 ;
        RECT 84.880 39.780 85.180 40.080 ;
        RECT 85.370 39.780 85.670 40.080 ;
        RECT 85.860 39.780 86.160 40.080 ;
        RECT 86.350 39.780 86.650 40.080 ;
        RECT 86.840 39.780 87.140 40.080 ;
        RECT 88.920 39.780 89.220 40.080 ;
        RECT 89.410 39.780 89.710 40.080 ;
        RECT 89.900 39.780 90.200 40.080 ;
        RECT 90.390 39.780 90.690 40.080 ;
        RECT 90.880 39.780 91.180 40.080 ;
        RECT 91.370 39.780 91.670 40.080 ;
        RECT 91.860 39.780 92.160 40.080 ;
        RECT 92.350 39.780 92.650 40.080 ;
        RECT 94.560 39.780 94.860 40.080 ;
        RECT 95.050 39.780 95.350 40.080 ;
        RECT 95.540 39.780 95.840 40.080 ;
        RECT 96.030 39.780 96.330 40.080 ;
        RECT 97.880 39.780 98.180 40.080 ;
        RECT 98.370 39.780 98.670 40.080 ;
        RECT 98.860 39.780 99.160 40.080 ;
        RECT 101.120 39.780 101.420 40.080 ;
        RECT 101.610 39.780 101.910 40.080 ;
        RECT 102.100 39.780 102.400 40.080 ;
        RECT 102.590 39.780 102.890 40.080 ;
        RECT 103.080 39.780 103.380 40.080 ;
        RECT 103.570 39.780 103.870 40.080 ;
        RECT 104.060 39.780 104.360 40.080 ;
        RECT 104.550 39.780 104.850 40.080 ;
        RECT 106.630 39.780 106.930 40.080 ;
        RECT 107.120 39.780 107.420 40.080 ;
        RECT 107.610 39.780 107.910 40.080 ;
        RECT 108.100 39.780 108.400 40.080 ;
        RECT 108.590 39.780 108.890 40.080 ;
        RECT 109.080 39.780 109.380 40.080 ;
        RECT 109.570 39.780 109.870 40.080 ;
        RECT 110.060 39.780 110.360 40.080 ;
        RECT 112.270 39.780 112.570 40.080 ;
        RECT 112.760 39.780 113.060 40.080 ;
        RECT 113.250 39.780 113.550 40.080 ;
        RECT 113.740 39.780 114.040 40.080 ;
        RECT 11.510 34.280 11.810 34.580 ;
        RECT 9.130 32.920 9.430 33.220 ;
        RECT 9.620 32.920 9.920 33.220 ;
        RECT 10.110 32.920 10.410 33.220 ;
        RECT 17.035 34.280 17.335 34.580 ;
        RECT 15.110 32.920 15.410 33.220 ;
        RECT 15.600 32.920 15.900 33.220 ;
        RECT 16.090 32.920 16.390 33.220 ;
        RECT 29.220 34.280 29.520 34.580 ;
        RECT 17.980 32.920 18.280 33.220 ;
        RECT 18.470 32.920 18.770 33.220 ;
        RECT 18.960 32.920 19.260 33.220 ;
        RECT 26.840 32.920 27.140 33.220 ;
        RECT 27.330 32.920 27.630 33.220 ;
        RECT 27.820 32.920 28.120 33.220 ;
        RECT 34.745 34.280 35.045 34.580 ;
        RECT 32.820 32.920 33.120 33.220 ;
        RECT 33.310 32.920 33.610 33.220 ;
        RECT 33.800 32.920 34.100 33.220 ;
        RECT 46.930 34.280 47.230 34.580 ;
        RECT 35.690 32.920 35.990 33.220 ;
        RECT 36.180 32.920 36.480 33.220 ;
        RECT 36.670 32.920 36.970 33.220 ;
        RECT 44.550 32.920 44.850 33.220 ;
        RECT 45.040 32.920 45.340 33.220 ;
        RECT 45.530 32.920 45.830 33.220 ;
        RECT 52.455 34.280 52.755 34.580 ;
        RECT 50.530 32.920 50.830 33.220 ;
        RECT 51.020 32.920 51.320 33.220 ;
        RECT 51.510 32.920 51.810 33.220 ;
        RECT 64.640 34.280 64.940 34.580 ;
        RECT 53.400 32.920 53.700 33.220 ;
        RECT 53.890 32.920 54.190 33.220 ;
        RECT 54.380 32.920 54.680 33.220 ;
        RECT 62.260 32.920 62.560 33.220 ;
        RECT 62.750 32.920 63.050 33.220 ;
        RECT 63.240 32.920 63.540 33.220 ;
        RECT 70.165 34.280 70.465 34.580 ;
        RECT 68.240 32.920 68.540 33.220 ;
        RECT 68.730 32.920 69.030 33.220 ;
        RECT 69.220 32.920 69.520 33.220 ;
        RECT 82.350 34.280 82.650 34.580 ;
        RECT 71.110 32.920 71.410 33.220 ;
        RECT 71.600 32.920 71.900 33.220 ;
        RECT 72.090 32.920 72.390 33.220 ;
        RECT 79.970 32.920 80.270 33.220 ;
        RECT 80.460 32.920 80.760 33.220 ;
        RECT 80.950 32.920 81.250 33.220 ;
        RECT 87.875 34.280 88.175 34.580 ;
        RECT 85.950 32.920 86.250 33.220 ;
        RECT 86.440 32.920 86.740 33.220 ;
        RECT 86.930 32.920 87.230 33.220 ;
        RECT 100.060 34.280 100.360 34.580 ;
        RECT 88.820 32.920 89.120 33.220 ;
        RECT 89.310 32.920 89.610 33.220 ;
        RECT 89.800 32.920 90.100 33.220 ;
        RECT 97.680 32.920 97.980 33.220 ;
        RECT 98.170 32.920 98.470 33.220 ;
        RECT 98.660 32.920 98.960 33.220 ;
        RECT 105.585 34.280 105.885 34.580 ;
        RECT 103.660 32.920 103.960 33.220 ;
        RECT 104.150 32.920 104.450 33.220 ;
        RECT 104.640 32.920 104.940 33.220 ;
        RECT 106.530 32.920 106.830 33.220 ;
        RECT 107.020 32.920 107.320 33.220 ;
        RECT 107.510 32.920 107.810 33.220 ;
      LAYER met1 ;
        RECT 22.390 48.590 26.660 48.950 ;
        RECT 31.240 48.590 32.740 48.950 ;
        RECT 40.100 48.590 44.370 48.950 ;
        RECT 48.950 48.590 50.450 48.950 ;
        RECT 57.810 48.590 62.080 48.950 ;
        RECT 66.660 48.590 68.160 48.950 ;
        RECT 75.520 48.590 79.790 48.950 ;
        RECT 84.370 48.590 85.870 48.950 ;
        RECT 93.230 48.590 97.500 48.950 ;
        RECT 102.080 48.590 103.580 48.950 ;
        RECT 23.005 47.590 23.365 48.590 ;
        RECT 31.790 47.590 32.150 48.590 ;
        RECT 40.715 47.590 41.075 48.590 ;
        RECT 49.500 47.590 49.860 48.590 ;
        RECT 58.425 47.590 58.785 48.590 ;
        RECT 67.210 47.590 67.570 48.590 ;
        RECT 76.135 47.590 76.495 48.590 ;
        RECT 84.920 47.590 85.280 48.590 ;
        RECT 93.845 47.590 94.205 48.590 ;
        RECT 102.630 47.590 102.990 48.590 ;
        RECT 14.620 47.230 23.365 47.590 ;
        RECT 24.315 47.230 41.075 47.590 ;
        RECT 42.025 47.230 58.785 47.590 ;
        RECT 59.735 47.230 76.495 47.590 ;
        RECT 77.445 47.230 94.205 47.590 ;
        RECT 95.155 47.230 106.360 47.590 ;
        RECT 14.620 42.000 14.980 47.230 ;
        RECT 6.350 41.640 14.980 42.000 ;
        RECT 15.980 41.670 105.050 42.150 ;
        RECT 106.000 42.000 106.360 47.230 ;
        RECT 109.500 44.500 110.500 45.515 ;
        RECT 106.000 41.640 115.500 42.000 ;
        RECT 6.350 34.610 6.710 41.640 ;
        RECT 7.500 39.690 114.280 40.170 ;
        RECT 115.140 34.610 115.500 41.640 ;
        RECT 6.350 34.250 17.395 34.610 ;
        RECT 18.345 34.250 35.105 34.610 ;
        RECT 36.055 34.250 52.815 34.610 ;
        RECT 53.765 34.250 70.525 34.610 ;
        RECT 71.475 34.250 88.235 34.610 ;
        RECT 89.185 34.250 105.945 34.610 ;
        RECT 106.895 34.250 115.500 34.610 ;
        RECT 9.560 33.250 9.920 34.250 ;
        RECT 18.345 33.250 18.705 34.250 ;
        RECT 27.270 33.250 27.630 34.250 ;
        RECT 36.055 33.250 36.415 34.250 ;
        RECT 44.980 33.250 45.340 34.250 ;
        RECT 53.765 33.250 54.125 34.250 ;
        RECT 62.690 33.250 63.050 34.250 ;
        RECT 71.475 33.250 71.835 34.250 ;
        RECT 80.400 33.250 80.760 34.250 ;
        RECT 89.185 33.250 89.545 34.250 ;
        RECT 98.110 33.250 98.470 34.250 ;
        RECT 106.895 33.250 107.255 34.250 ;
        RECT 8.970 32.890 10.470 33.250 ;
        RECT 15.050 32.890 19.320 33.250 ;
        RECT 26.680 32.890 28.180 33.250 ;
        RECT 32.760 32.890 37.030 33.250 ;
        RECT 44.390 32.890 45.890 33.250 ;
        RECT 50.470 32.890 54.740 33.250 ;
        RECT 62.100 32.890 63.600 33.250 ;
        RECT 68.180 32.890 72.450 33.250 ;
        RECT 79.810 32.890 81.310 33.250 ;
        RECT 85.890 32.890 90.160 33.250 ;
        RECT 97.520 32.890 99.020 33.250 ;
        RECT 103.600 32.890 107.870 33.250 ;
      LAYER via ;
        RECT 19.500 41.770 19.760 42.030 ;
        RECT 19.870 41.770 20.130 42.030 ;
        RECT 20.240 41.770 20.500 42.030 ;
        RECT 25.500 41.770 25.760 42.030 ;
        RECT 25.870 41.770 26.130 42.030 ;
        RECT 26.240 41.770 26.500 42.030 ;
        RECT 31.500 41.770 31.760 42.030 ;
        RECT 31.870 41.770 32.130 42.030 ;
        RECT 32.240 41.770 32.500 42.030 ;
        RECT 37.500 41.770 37.760 42.030 ;
        RECT 37.870 41.770 38.130 42.030 ;
        RECT 38.240 41.770 38.500 42.030 ;
        RECT 43.500 41.770 43.760 42.030 ;
        RECT 43.870 41.770 44.130 42.030 ;
        RECT 44.240 41.770 44.500 42.030 ;
        RECT 49.500 41.770 49.760 42.030 ;
        RECT 49.870 41.770 50.130 42.030 ;
        RECT 50.240 41.770 50.500 42.030 ;
        RECT 55.500 41.770 55.760 42.030 ;
        RECT 55.870 41.770 56.130 42.030 ;
        RECT 56.240 41.770 56.500 42.030 ;
        RECT 61.500 41.770 61.760 42.030 ;
        RECT 61.870 41.770 62.130 42.030 ;
        RECT 62.240 41.770 62.500 42.030 ;
        RECT 67.500 41.770 67.760 42.030 ;
        RECT 67.870 41.770 68.130 42.030 ;
        RECT 68.240 41.770 68.500 42.030 ;
        RECT 73.500 41.770 73.760 42.030 ;
        RECT 73.870 41.770 74.130 42.030 ;
        RECT 74.240 41.770 74.500 42.030 ;
        RECT 79.500 41.770 79.760 42.030 ;
        RECT 79.870 41.770 80.130 42.030 ;
        RECT 80.240 41.770 80.500 42.030 ;
        RECT 85.500 41.770 85.760 42.030 ;
        RECT 85.870 41.770 86.130 42.030 ;
        RECT 86.240 41.770 86.500 42.030 ;
        RECT 91.500 41.770 91.760 42.030 ;
        RECT 91.870 41.770 92.130 42.030 ;
        RECT 92.240 41.770 92.500 42.030 ;
        RECT 97.500 41.770 97.760 42.030 ;
        RECT 97.870 41.770 98.130 42.030 ;
        RECT 98.240 41.770 98.500 42.030 ;
        RECT 103.500 41.770 103.760 42.030 ;
        RECT 103.870 41.770 104.130 42.030 ;
        RECT 104.240 41.770 104.500 42.030 ;
        RECT 109.570 45.100 109.910 45.440 ;
        RECT 110.090 45.100 110.430 45.440 ;
        RECT 109.570 44.580 109.910 44.920 ;
        RECT 110.090 44.580 110.430 44.920 ;
        RECT 7.500 39.790 7.760 40.050 ;
        RECT 7.870 39.790 8.130 40.050 ;
        RECT 8.240 39.790 8.500 40.050 ;
        RECT 13.500 39.790 13.760 40.050 ;
        RECT 13.870 39.790 14.130 40.050 ;
        RECT 14.240 39.790 14.500 40.050 ;
        RECT 19.500 39.790 19.760 40.050 ;
        RECT 19.870 39.790 20.130 40.050 ;
        RECT 20.240 39.790 20.500 40.050 ;
        RECT 25.500 39.790 25.760 40.050 ;
        RECT 25.870 39.790 26.130 40.050 ;
        RECT 26.240 39.790 26.500 40.050 ;
        RECT 31.500 39.790 31.760 40.050 ;
        RECT 31.870 39.790 32.130 40.050 ;
        RECT 32.240 39.790 32.500 40.050 ;
        RECT 37.500 39.790 37.760 40.050 ;
        RECT 37.870 39.790 38.130 40.050 ;
        RECT 38.240 39.790 38.500 40.050 ;
        RECT 43.500 39.790 43.760 40.050 ;
        RECT 43.870 39.790 44.130 40.050 ;
        RECT 44.240 39.790 44.500 40.050 ;
        RECT 49.500 39.790 49.760 40.050 ;
        RECT 49.870 39.790 50.130 40.050 ;
        RECT 50.240 39.790 50.500 40.050 ;
        RECT 55.500 39.790 55.760 40.050 ;
        RECT 55.870 39.790 56.130 40.050 ;
        RECT 56.240 39.790 56.500 40.050 ;
        RECT 61.500 39.790 61.760 40.050 ;
        RECT 61.870 39.790 62.130 40.050 ;
        RECT 62.240 39.790 62.500 40.050 ;
        RECT 67.500 39.790 67.760 40.050 ;
        RECT 67.870 39.790 68.130 40.050 ;
        RECT 68.240 39.790 68.500 40.050 ;
        RECT 73.500 39.790 73.760 40.050 ;
        RECT 73.870 39.790 74.130 40.050 ;
        RECT 74.240 39.790 74.500 40.050 ;
        RECT 79.500 39.790 79.760 40.050 ;
        RECT 79.870 39.790 80.130 40.050 ;
        RECT 80.240 39.790 80.500 40.050 ;
        RECT 85.500 39.790 85.760 40.050 ;
        RECT 85.870 39.790 86.130 40.050 ;
        RECT 86.240 39.790 86.500 40.050 ;
        RECT 91.500 39.790 91.760 40.050 ;
        RECT 91.870 39.790 92.130 40.050 ;
        RECT 92.240 39.790 92.500 40.050 ;
        RECT 97.500 39.790 97.760 40.050 ;
        RECT 97.870 39.790 98.130 40.050 ;
        RECT 98.240 39.790 98.500 40.050 ;
        RECT 103.500 39.790 103.760 40.050 ;
        RECT 103.870 39.790 104.130 40.050 ;
        RECT 104.240 39.790 104.500 40.050 ;
        RECT 109.500 39.790 109.760 40.050 ;
        RECT 109.870 39.790 110.130 40.050 ;
        RECT 110.240 39.790 110.500 40.050 ;
        RECT 113.280 39.790 113.540 40.050 ;
        RECT 113.650 39.790 113.910 40.050 ;
        RECT 114.020 39.790 114.280 40.050 ;
      LAYER met2 ;
        RECT 109.500 44.500 110.500 45.515 ;
        RECT 19.500 41.700 20.500 42.100 ;
        RECT 25.500 41.700 26.500 42.100 ;
        RECT 31.500 41.700 32.500 42.100 ;
        RECT 37.500 41.700 38.500 42.100 ;
        RECT 43.500 41.700 44.500 42.100 ;
        RECT 49.500 41.700 50.500 42.100 ;
        RECT 55.500 41.700 56.500 42.100 ;
        RECT 61.500 41.700 62.500 42.100 ;
        RECT 67.500 41.700 68.500 42.100 ;
        RECT 73.500 41.700 74.500 42.100 ;
        RECT 79.500 41.700 80.500 42.100 ;
        RECT 85.500 41.700 86.500 42.100 ;
        RECT 91.500 41.700 92.500 42.100 ;
        RECT 97.500 41.700 98.500 42.100 ;
        RECT 103.500 41.700 104.500 42.100 ;
        RECT 7.500 39.720 8.500 40.120 ;
        RECT 13.500 39.720 14.500 40.120 ;
        RECT 19.500 39.720 20.500 40.120 ;
        RECT 25.500 39.720 26.500 40.120 ;
        RECT 31.500 39.720 32.500 40.120 ;
        RECT 37.500 39.720 38.500 40.120 ;
        RECT 43.500 39.720 44.500 40.120 ;
        RECT 49.500 39.720 50.500 40.120 ;
        RECT 55.500 39.720 56.500 40.120 ;
        RECT 61.500 39.720 62.500 40.120 ;
        RECT 67.500 39.720 68.500 40.120 ;
        RECT 73.500 39.720 74.500 40.120 ;
        RECT 79.500 39.720 80.500 40.120 ;
        RECT 85.500 39.720 86.500 40.120 ;
        RECT 91.500 39.720 92.500 40.120 ;
        RECT 97.500 39.720 98.500 40.120 ;
        RECT 103.500 39.720 104.500 40.120 ;
        RECT 109.500 39.720 110.500 40.120 ;
        RECT 113.280 39.720 114.280 40.120 ;
      LAYER via2 ;
        RECT 109.540 45.070 109.940 45.470 ;
        RECT 110.060 45.070 110.460 45.470 ;
        RECT 109.540 44.550 109.940 44.950 ;
        RECT 110.060 44.550 110.460 44.950 ;
        RECT 19.600 41.750 19.900 42.050 ;
        RECT 20.100 41.750 20.400 42.050 ;
        RECT 25.600 41.750 25.900 42.050 ;
        RECT 26.100 41.750 26.400 42.050 ;
        RECT 31.600 41.750 31.900 42.050 ;
        RECT 32.100 41.750 32.400 42.050 ;
        RECT 37.600 41.750 37.900 42.050 ;
        RECT 38.100 41.750 38.400 42.050 ;
        RECT 43.600 41.750 43.900 42.050 ;
        RECT 44.100 41.750 44.400 42.050 ;
        RECT 49.600 41.750 49.900 42.050 ;
        RECT 50.100 41.750 50.400 42.050 ;
        RECT 55.600 41.750 55.900 42.050 ;
        RECT 56.100 41.750 56.400 42.050 ;
        RECT 61.600 41.750 61.900 42.050 ;
        RECT 62.100 41.750 62.400 42.050 ;
        RECT 67.600 41.750 67.900 42.050 ;
        RECT 68.100 41.750 68.400 42.050 ;
        RECT 73.600 41.750 73.900 42.050 ;
        RECT 74.100 41.750 74.400 42.050 ;
        RECT 79.600 41.750 79.900 42.050 ;
        RECT 80.100 41.750 80.400 42.050 ;
        RECT 85.600 41.750 85.900 42.050 ;
        RECT 86.100 41.750 86.400 42.050 ;
        RECT 91.600 41.750 91.900 42.050 ;
        RECT 92.100 41.750 92.400 42.050 ;
        RECT 97.600 41.750 97.900 42.050 ;
        RECT 98.100 41.750 98.400 42.050 ;
        RECT 103.600 41.750 103.900 42.050 ;
        RECT 104.100 41.750 104.400 42.050 ;
        RECT 7.600 39.770 7.900 40.070 ;
        RECT 8.100 39.770 8.400 40.070 ;
        RECT 13.600 39.770 13.900 40.070 ;
        RECT 14.100 39.770 14.400 40.070 ;
        RECT 19.600 39.770 19.900 40.070 ;
        RECT 20.100 39.770 20.400 40.070 ;
        RECT 25.600 39.770 25.900 40.070 ;
        RECT 26.100 39.770 26.400 40.070 ;
        RECT 31.600 39.770 31.900 40.070 ;
        RECT 32.100 39.770 32.400 40.070 ;
        RECT 37.600 39.770 37.900 40.070 ;
        RECT 38.100 39.770 38.400 40.070 ;
        RECT 43.600 39.770 43.900 40.070 ;
        RECT 44.100 39.770 44.400 40.070 ;
        RECT 49.600 39.770 49.900 40.070 ;
        RECT 50.100 39.770 50.400 40.070 ;
        RECT 55.600 39.770 55.900 40.070 ;
        RECT 56.100 39.770 56.400 40.070 ;
        RECT 61.600 39.770 61.900 40.070 ;
        RECT 62.100 39.770 62.400 40.070 ;
        RECT 67.600 39.770 67.900 40.070 ;
        RECT 68.100 39.770 68.400 40.070 ;
        RECT 73.600 39.770 73.900 40.070 ;
        RECT 74.100 39.770 74.400 40.070 ;
        RECT 79.600 39.770 79.900 40.070 ;
        RECT 80.100 39.770 80.400 40.070 ;
        RECT 85.600 39.770 85.900 40.070 ;
        RECT 86.100 39.770 86.400 40.070 ;
        RECT 91.600 39.770 91.900 40.070 ;
        RECT 92.100 39.770 92.400 40.070 ;
        RECT 97.600 39.770 97.900 40.070 ;
        RECT 98.100 39.770 98.400 40.070 ;
        RECT 103.600 39.770 103.900 40.070 ;
        RECT 104.100 39.770 104.400 40.070 ;
        RECT 109.600 39.770 109.900 40.070 ;
        RECT 110.100 39.770 110.400 40.070 ;
        RECT 113.380 39.770 113.680 40.070 ;
        RECT 113.880 39.770 114.180 40.070 ;
      LAYER met3 ;
        RECT 19.500 41.670 20.500 42.150 ;
        RECT 25.500 41.670 26.500 42.150 ;
        RECT 31.500 41.670 32.500 42.150 ;
        RECT 37.500 41.670 38.500 42.150 ;
        RECT 43.500 41.670 44.500 42.150 ;
        RECT 49.500 41.670 50.500 42.150 ;
        RECT 55.500 41.670 56.500 42.150 ;
        RECT 61.500 41.670 62.500 42.150 ;
        RECT 67.500 41.670 68.500 42.150 ;
        RECT 73.500 41.670 74.500 42.150 ;
        RECT 79.500 41.670 80.500 42.150 ;
        RECT 85.500 41.670 86.500 42.150 ;
        RECT 91.500 41.670 92.500 42.150 ;
        RECT 97.500 41.670 98.500 42.150 ;
        RECT 103.500 41.670 104.500 42.150 ;
        RECT 109.500 41.670 110.500 45.515 ;
        RECT 7.500 40.170 114.280 41.670 ;
        RECT 7.500 39.690 8.500 40.170 ;
        RECT 13.500 39.690 14.500 40.170 ;
        RECT 19.500 39.690 20.500 40.170 ;
        RECT 25.500 39.690 26.500 40.170 ;
        RECT 31.500 39.690 32.500 40.170 ;
        RECT 37.500 39.690 38.500 40.170 ;
        RECT 43.500 39.690 44.500 40.170 ;
        RECT 49.500 39.690 50.500 40.170 ;
        RECT 55.500 39.690 56.500 40.170 ;
        RECT 61.500 39.690 62.500 40.170 ;
        RECT 67.500 39.690 68.500 40.170 ;
        RECT 73.500 39.690 74.500 40.170 ;
        RECT 79.500 39.690 80.500 40.170 ;
        RECT 85.500 39.690 86.500 40.170 ;
        RECT 91.500 39.690 92.500 40.170 ;
        RECT 97.500 39.690 98.500 40.170 ;
        RECT 103.500 39.690 104.500 40.170 ;
        RECT 109.500 39.690 110.500 40.170 ;
        RECT 113.280 39.690 114.280 40.170 ;
  END
END vco_w6_r100
END LIBRARY

