magic
tech sky130A
magscale 1 2
timestamp 1623172581
<< ndiff >>
rect 1054 11992 1082 12024
<< pdiff >>
rect 1052 12300 1084 12334
<< psubdiff >>
rect 21698 6000 21700 6100
rect 21800 6000 21900 6100
rect 22000 6000 22098 6100
<< locali >>
rect 1327 12275 1496 12335
rect 781 12099 873 12245
rect 1786 12216 1830 12260
rect 954 12118 978 12144
rect 21698 6000 21700 6100
rect 21800 6080 21900 6100
rect 22000 6080 22098 6100
rect 21800 6020 21818 6080
rect 21878 6020 21900 6080
rect 22000 6020 22018 6080
rect 22078 6020 22098 6080
rect 21800 6000 21900 6020
rect 22000 6000 22098 6020
<< viali >>
rect 7318 14420 7378 14480
rect 7418 14420 7478 14480
rect 7518 14420 7578 14480
rect 7618 14420 7678 14480
rect 14518 14420 14578 14480
rect 14618 14420 14678 14480
rect 14718 14420 14778 14480
rect 14818 14420 14878 14480
rect 21718 14420 21778 14480
rect 21818 14420 21878 14480
rect 21918 14420 21978 14480
rect 22018 14420 22078 14480
rect 28918 14420 28978 14480
rect 29018 14420 29078 14480
rect 29118 14420 29178 14480
rect 29218 14420 29278 14480
rect 7318 6020 7378 6080
rect 7418 6020 7478 6080
rect 7518 6020 7578 6080
rect 7618 6020 7678 6080
rect 14518 6020 14578 6080
rect 14618 6020 14678 6080
rect 14718 6020 14778 6080
rect 14818 6020 14878 6080
rect 21718 6020 21778 6080
rect 21818 6020 21878 6080
rect 21918 6020 21978 6080
rect 22018 6020 22078 6080
rect 28918 6020 28978 6080
rect 29018 6020 29078 6080
rect 29118 6020 29178 6080
rect 29218 6020 29278 6080
<< metal1 >>
rect 7298 14480 7698 14500
rect 7298 14420 7318 14480
rect 7384 14420 7396 14480
rect 7600 14420 7612 14480
rect 7678 14420 7698 14480
rect 7298 14400 7698 14420
rect 14498 14480 14898 14500
rect 14498 14420 14518 14480
rect 14584 14420 14596 14480
rect 14800 14420 14812 14480
rect 14878 14420 14898 14480
rect 14498 14400 14898 14420
rect 21698 14480 22098 14500
rect 21698 14420 21718 14480
rect 21784 14420 21796 14480
rect 22000 14420 22012 14480
rect 22078 14420 22098 14480
rect 21698 14400 22098 14420
rect 28898 14480 29298 14500
rect 28898 14420 28918 14480
rect 28984 14420 28996 14480
rect 29200 14420 29212 14480
rect 29278 14420 29298 14480
rect 28898 14400 29298 14420
rect 3200 13562 4072 13580
rect 3200 13502 3724 13562
rect 3784 13502 3796 13562
rect 3856 13502 3868 13562
rect 3928 13502 3940 13562
rect 4000 13502 4012 13562
rect 3200 13484 4072 13502
rect 10924 13562 11272 13580
rect 10984 13502 10996 13562
rect 11056 13502 11068 13562
rect 11128 13502 11140 13562
rect 11200 13502 11212 13562
rect 10924 13484 11272 13502
rect 18124 13562 18472 13580
rect 18184 13502 18196 13562
rect 18256 13502 18268 13562
rect 18328 13502 18340 13562
rect 18400 13502 18412 13562
rect 18124 13484 18472 13502
rect 25324 13562 25672 13580
rect 25384 13502 25396 13562
rect 25456 13502 25468 13562
rect 25528 13502 25540 13562
rect 25600 13502 25612 13562
rect 25324 13484 25672 13502
rect 32524 13562 32872 13580
rect 32584 13502 32596 13562
rect 32656 13502 32668 13562
rect 32728 13502 32740 13562
rect 32800 13502 32812 13562
rect 32524 13484 32872 13502
rect 9336 12652 9634 12780
rect 15248 12654 15546 12782
rect 21152 12652 21450 12780
rect 27044 12652 27342 12780
rect 2950 12474 4098 12492
rect 2950 12414 3724 12474
rect 3784 12414 3796 12474
rect 3856 12414 3868 12474
rect 3928 12414 3940 12474
rect 4000 12414 4012 12474
rect 4072 12414 4098 12474
rect 2950 12396 4098 12414
rect 98 11930 498 11948
rect 98 11870 124 11930
rect 184 11870 196 11930
rect 256 11870 268 11930
rect 328 11870 340 11930
rect 400 11870 412 11930
rect 472 11870 498 11930
rect 98 11852 498 11870
rect 3002 11386 4072 11404
rect 3002 11326 3724 11386
rect 3784 11326 3796 11386
rect 3856 11326 3868 11386
rect 3928 11326 3940 11386
rect 4000 11326 4012 11386
rect 3002 11308 4072 11326
rect 10924 11386 11272 11404
rect 10984 11326 10996 11386
rect 11056 11326 11068 11386
rect 11128 11326 11140 11386
rect 11200 11326 11212 11386
rect 10924 11308 11272 11326
rect 18124 11386 18472 11404
rect 18184 11326 18196 11386
rect 18256 11326 18268 11386
rect 18328 11326 18340 11386
rect 18400 11326 18412 11386
rect 18124 11308 18472 11326
rect 25324 11386 25672 11404
rect 25384 11326 25396 11386
rect 25456 11326 25468 11386
rect 25528 11326 25540 11386
rect 25600 11326 25612 11386
rect 25324 11308 25672 11326
rect 32524 11385 34290 11404
rect 32584 11325 32596 11385
rect 32656 11325 32668 11385
rect 32728 11325 32740 11385
rect 32800 11325 32812 11385
rect 32872 11325 34290 11385
rect 32524 11308 34290 11325
rect 32498 11307 32898 11308
rect 31002 10762 31520 10860
rect 0 9210 4072 9228
rect 0 9150 3724 9210
rect 3784 9150 3796 9210
rect 3856 9150 3868 9210
rect 3928 9150 3940 9210
rect 4000 9150 4012 9210
rect 0 9132 4072 9150
rect 10924 9210 11272 9228
rect 10984 9150 10996 9210
rect 11056 9150 11068 9210
rect 11128 9150 11140 9210
rect 11200 9150 11212 9210
rect 10924 9132 11272 9150
rect 18124 9210 18472 9228
rect 18184 9150 18196 9210
rect 18256 9150 18268 9210
rect 18328 9150 18340 9210
rect 18400 9150 18412 9210
rect 18124 9132 18472 9150
rect 25324 9210 25672 9228
rect 25384 9150 25396 9210
rect 25456 9150 25468 9210
rect 25528 9150 25540 9210
rect 25600 9150 25612 9210
rect 25324 9132 25672 9150
rect 32524 9210 35889 9228
rect 32584 9150 32596 9210
rect 32656 9150 32668 9210
rect 32728 9150 32740 9210
rect 32800 9150 32812 9210
rect 32872 9150 35889 9210
rect 32524 9132 35889 9150
rect 6144 7756 6442 7884
rect 12044 7754 12342 7882
rect 17956 7754 18254 7882
rect 23852 7754 24150 7882
rect 29768 7754 30066 7882
rect 0 7034 4072 7052
rect 0 6974 3724 7034
rect 3784 6974 3796 7034
rect 3856 6974 3868 7034
rect 3928 6974 3940 7034
rect 4000 6974 4012 7034
rect 0 6956 4072 6974
rect 10924 7034 11272 7052
rect 10984 6974 10996 7034
rect 11056 6974 11068 7034
rect 11128 6974 11140 7034
rect 11200 6974 11212 7034
rect 10924 6956 11272 6974
rect 25324 7034 25672 7052
rect 25384 6974 25396 7034
rect 25456 6974 25468 7034
rect 25528 6974 25540 7034
rect 25600 6974 25612 7034
rect 25324 6956 25672 6974
rect 32524 7034 35888 7052
rect 32584 6974 32596 7034
rect 32656 6974 32668 7034
rect 32728 6974 32740 7034
rect 32800 6974 32812 7034
rect 32872 6974 35888 7034
rect 32524 6956 35888 6974
rect 7298 6080 7698 6100
rect 7298 6020 7318 6080
rect 7384 6020 7396 6080
rect 7600 6020 7612 6080
rect 7678 6020 7698 6080
rect 7298 6000 7698 6020
rect 14498 6080 14898 6100
rect 14498 6020 14518 6080
rect 14584 6020 14596 6080
rect 14800 6020 14812 6080
rect 14878 6020 14898 6080
rect 14498 6000 14898 6020
rect 21698 6080 22098 6100
rect 21698 6020 21718 6080
rect 21784 6020 21796 6080
rect 22000 6020 22012 6080
rect 22078 6020 22098 6080
rect 21698 6000 22098 6020
rect 28898 6080 29298 6100
rect 28898 6020 28918 6080
rect 28984 6020 28996 6080
rect 29200 6020 29212 6080
rect 29278 6020 29298 6080
rect 28898 6000 29298 6020
<< via1 >>
rect 7324 14420 7378 14480
rect 7378 14420 7384 14480
rect 7396 14420 7418 14480
rect 7418 14420 7456 14480
rect 7468 14420 7478 14480
rect 7478 14420 7518 14480
rect 7518 14420 7528 14480
rect 7540 14420 7578 14480
rect 7578 14420 7600 14480
rect 7612 14420 7618 14480
rect 7618 14420 7672 14480
rect 14524 14420 14578 14480
rect 14578 14420 14584 14480
rect 14596 14420 14618 14480
rect 14618 14420 14656 14480
rect 14668 14420 14678 14480
rect 14678 14420 14718 14480
rect 14718 14420 14728 14480
rect 14740 14420 14778 14480
rect 14778 14420 14800 14480
rect 14812 14420 14818 14480
rect 14818 14420 14872 14480
rect 21724 14420 21778 14480
rect 21778 14420 21784 14480
rect 21796 14420 21818 14480
rect 21818 14420 21856 14480
rect 21868 14420 21878 14480
rect 21878 14420 21918 14480
rect 21918 14420 21928 14480
rect 21940 14420 21978 14480
rect 21978 14420 22000 14480
rect 22012 14420 22018 14480
rect 22018 14420 22072 14480
rect 28924 14420 28978 14480
rect 28978 14420 28984 14480
rect 28996 14420 29018 14480
rect 29018 14420 29056 14480
rect 29068 14420 29078 14480
rect 29078 14420 29118 14480
rect 29118 14420 29128 14480
rect 29140 14420 29178 14480
rect 29178 14420 29200 14480
rect 29212 14420 29218 14480
rect 29218 14420 29272 14480
rect 3724 13502 3784 13562
rect 3796 13502 3856 13562
rect 3868 13502 3928 13562
rect 3940 13502 4000 13562
rect 4012 13502 4072 13562
rect 10924 13502 10984 13562
rect 10996 13502 11056 13562
rect 11068 13502 11128 13562
rect 11140 13502 11200 13562
rect 11212 13502 11272 13562
rect 18124 13502 18184 13562
rect 18196 13502 18256 13562
rect 18268 13502 18328 13562
rect 18340 13502 18400 13562
rect 18412 13502 18472 13562
rect 25324 13502 25384 13562
rect 25396 13502 25456 13562
rect 25468 13502 25528 13562
rect 25540 13502 25600 13562
rect 25612 13502 25672 13562
rect 32524 13502 32584 13562
rect 32596 13502 32656 13562
rect 32668 13502 32728 13562
rect 32740 13502 32800 13562
rect 32812 13502 32872 13562
rect 3724 12414 3784 12474
rect 3796 12414 3856 12474
rect 3868 12414 3928 12474
rect 3940 12414 4000 12474
rect 4012 12414 4072 12474
rect 124 11870 184 11930
rect 196 11870 256 11930
rect 268 11870 328 11930
rect 340 11870 400 11930
rect 412 11870 472 11930
rect 3724 11326 3784 11386
rect 3796 11326 3856 11386
rect 3868 11326 3928 11386
rect 3940 11326 4000 11386
rect 4012 11326 4072 11386
rect 10924 11326 10984 11386
rect 10996 11326 11056 11386
rect 11068 11326 11128 11386
rect 11140 11326 11200 11386
rect 11212 11326 11272 11386
rect 18124 11326 18184 11386
rect 18196 11326 18256 11386
rect 18268 11326 18328 11386
rect 18340 11326 18400 11386
rect 18412 11326 18472 11386
rect 25324 11326 25384 11386
rect 25396 11326 25456 11386
rect 25468 11326 25528 11386
rect 25540 11326 25600 11386
rect 25612 11326 25672 11386
rect 32524 11325 32584 11385
rect 32596 11325 32656 11385
rect 32668 11325 32728 11385
rect 32740 11325 32800 11385
rect 32812 11325 32872 11385
rect 3724 9150 3784 9210
rect 3796 9150 3856 9210
rect 3868 9150 3928 9210
rect 3940 9150 4000 9210
rect 4012 9150 4072 9210
rect 10924 9150 10984 9210
rect 10996 9150 11056 9210
rect 11068 9150 11128 9210
rect 11140 9150 11200 9210
rect 11212 9150 11272 9210
rect 18124 9150 18184 9210
rect 18196 9150 18256 9210
rect 18268 9150 18328 9210
rect 18340 9150 18400 9210
rect 18412 9150 18472 9210
rect 25324 9150 25384 9210
rect 25396 9150 25456 9210
rect 25468 9150 25528 9210
rect 25540 9150 25600 9210
rect 25612 9150 25672 9210
rect 32524 9150 32584 9210
rect 32596 9150 32656 9210
rect 32668 9150 32728 9210
rect 32740 9150 32800 9210
rect 32812 9150 32872 9210
rect 3724 6974 3784 7034
rect 3796 6974 3856 7034
rect 3868 6974 3928 7034
rect 3940 6974 4000 7034
rect 4012 6974 4072 7034
rect 10924 6974 10984 7034
rect 10996 6974 11056 7034
rect 11068 6974 11128 7034
rect 11140 6974 11200 7034
rect 11212 6974 11272 7034
rect 25324 6974 25384 7034
rect 25396 6974 25456 7034
rect 25468 6974 25528 7034
rect 25540 6974 25600 7034
rect 25612 6974 25672 7034
rect 32524 6974 32584 7034
rect 32596 6974 32656 7034
rect 32668 6974 32728 7034
rect 32740 6974 32800 7034
rect 32812 6974 32872 7034
rect 7324 6020 7378 6080
rect 7378 6020 7384 6080
rect 7396 6020 7418 6080
rect 7418 6020 7456 6080
rect 7468 6020 7478 6080
rect 7478 6020 7518 6080
rect 7518 6020 7528 6080
rect 7540 6020 7578 6080
rect 7578 6020 7600 6080
rect 7612 6020 7618 6080
rect 7618 6020 7672 6080
rect 14524 6020 14578 6080
rect 14578 6020 14584 6080
rect 14596 6020 14618 6080
rect 14618 6020 14656 6080
rect 14668 6020 14678 6080
rect 14678 6020 14718 6080
rect 14718 6020 14728 6080
rect 14740 6020 14778 6080
rect 14778 6020 14800 6080
rect 14812 6020 14818 6080
rect 14818 6020 14872 6080
rect 21724 6020 21778 6080
rect 21778 6020 21784 6080
rect 21796 6020 21818 6080
rect 21818 6020 21856 6080
rect 21868 6020 21878 6080
rect 21878 6020 21918 6080
rect 21918 6020 21928 6080
rect 21940 6020 21978 6080
rect 21978 6020 22000 6080
rect 22012 6020 22018 6080
rect 22018 6020 22072 6080
rect 28924 6020 28978 6080
rect 28978 6020 28984 6080
rect 28996 6020 29018 6080
rect 29018 6020 29056 6080
rect 29068 6020 29078 6080
rect 29078 6020 29118 6080
rect 29118 6020 29128 6080
rect 29140 6020 29178 6080
rect 29178 6020 29200 6080
rect 29212 6020 29218 6080
rect 29218 6020 29272 6080
<< metal2 >>
rect 7298 14482 7698 14500
rect 7298 14480 7334 14482
rect 7398 14480 7422 14482
rect 7486 14480 7510 14482
rect 7574 14480 7598 14482
rect 7662 14480 7698 14482
rect 7298 14420 7324 14480
rect 7672 14420 7698 14480
rect 7298 14418 7334 14420
rect 7398 14418 7422 14420
rect 7486 14418 7510 14420
rect 7574 14418 7598 14420
rect 7662 14418 7698 14420
rect 7298 14400 7698 14418
rect 14498 14482 14898 14500
rect 14498 14480 14534 14482
rect 14598 14480 14622 14482
rect 14686 14480 14710 14482
rect 14774 14480 14798 14482
rect 14862 14480 14898 14482
rect 14498 14420 14524 14480
rect 14872 14420 14898 14480
rect 14498 14418 14534 14420
rect 14598 14418 14622 14420
rect 14686 14418 14710 14420
rect 14774 14418 14798 14420
rect 14862 14418 14898 14420
rect 14498 14400 14898 14418
rect 21698 14482 22098 14500
rect 21698 14480 21734 14482
rect 21798 14480 21822 14482
rect 21886 14480 21910 14482
rect 21974 14480 21998 14482
rect 22062 14480 22098 14482
rect 21698 14420 21724 14480
rect 22072 14420 22098 14480
rect 21698 14418 21734 14420
rect 21798 14418 21822 14420
rect 21886 14418 21910 14420
rect 21974 14418 21998 14420
rect 22062 14418 22098 14420
rect 21698 14400 22098 14418
rect 28898 14482 29298 14500
rect 28898 14480 28934 14482
rect 28998 14480 29022 14482
rect 29086 14480 29110 14482
rect 29174 14480 29198 14482
rect 29262 14480 29298 14482
rect 28898 14420 28924 14480
rect 29272 14420 29298 14480
rect 28898 14418 28934 14420
rect 28998 14418 29022 14420
rect 29086 14418 29110 14420
rect 29174 14418 29198 14420
rect 29262 14418 29298 14420
rect 28898 14400 29298 14418
rect 9364 14134 9524 14334
rect 15264 14134 15424 14334
rect 21164 14134 21324 14334
rect 27064 14134 27224 14334
rect 3698 13564 4098 13580
rect 3698 13562 3734 13564
rect 3798 13562 3822 13564
rect 3886 13562 3910 13564
rect 3974 13562 3998 13564
rect 4062 13562 4098 13564
rect 3698 13502 3724 13562
rect 4072 13502 4098 13562
rect 3698 13500 3734 13502
rect 3798 13500 3822 13502
rect 3886 13500 3910 13502
rect 3974 13500 3998 13502
rect 4062 13500 4098 13502
rect 3698 13484 4098 13500
rect 10898 13564 11298 13580
rect 10898 13562 10934 13564
rect 10998 13562 11022 13564
rect 11086 13562 11110 13564
rect 11174 13562 11198 13564
rect 11262 13562 11298 13564
rect 10898 13502 10924 13562
rect 11272 13502 11298 13562
rect 10898 13500 10934 13502
rect 10998 13500 11022 13502
rect 11086 13500 11110 13502
rect 11174 13500 11198 13502
rect 11262 13500 11298 13502
rect 10898 13484 11298 13500
rect 18098 13564 18498 13580
rect 18098 13562 18134 13564
rect 18198 13562 18222 13564
rect 18286 13562 18310 13564
rect 18374 13562 18398 13564
rect 18462 13562 18498 13564
rect 18098 13502 18124 13562
rect 18472 13502 18498 13562
rect 18098 13500 18134 13502
rect 18198 13500 18222 13502
rect 18286 13500 18310 13502
rect 18374 13500 18398 13502
rect 18462 13500 18498 13502
rect 18098 13484 18498 13500
rect 25298 13564 25698 13580
rect 25298 13562 25334 13564
rect 25398 13562 25422 13564
rect 25486 13562 25510 13564
rect 25574 13562 25598 13564
rect 25662 13562 25698 13564
rect 25298 13502 25324 13562
rect 25672 13502 25698 13562
rect 25298 13500 25334 13502
rect 25398 13500 25422 13502
rect 25486 13500 25510 13502
rect 25574 13500 25598 13502
rect 25662 13500 25698 13502
rect 25298 13484 25698 13500
rect 32498 13564 32898 13580
rect 32498 13562 32534 13564
rect 32598 13562 32622 13564
rect 32686 13562 32710 13564
rect 32774 13562 32798 13564
rect 32862 13562 32898 13564
rect 32498 13502 32524 13562
rect 32872 13502 32898 13562
rect 32498 13500 32534 13502
rect 32598 13500 32622 13502
rect 32686 13500 32710 13502
rect 32774 13500 32798 13502
rect 32862 13500 32898 13502
rect 32498 13484 32898 13500
rect 3698 12476 4098 12492
rect 3698 12474 3734 12476
rect 3798 12474 3822 12476
rect 3886 12474 3910 12476
rect 3974 12474 3998 12476
rect 4062 12474 4098 12476
rect 3698 12414 3724 12474
rect 4072 12414 4098 12474
rect 3698 12412 3734 12414
rect 3798 12412 3822 12414
rect 3886 12412 3910 12414
rect 3974 12412 3998 12414
rect 4062 12412 4098 12414
rect 3698 12396 4098 12412
rect 98 11932 498 11948
rect 98 11930 134 11932
rect 198 11930 222 11932
rect 286 11930 310 11932
rect 374 11930 398 11932
rect 462 11930 498 11932
rect 98 11870 124 11930
rect 472 11870 498 11930
rect 98 11868 134 11870
rect 198 11868 222 11870
rect 286 11868 310 11870
rect 374 11868 398 11870
rect 462 11868 498 11870
rect 98 11852 498 11868
rect 3698 11388 4098 11404
rect 3698 11386 3734 11388
rect 3798 11386 3822 11388
rect 3886 11386 3910 11388
rect 3974 11386 3998 11388
rect 4062 11386 4098 11388
rect 3698 11326 3724 11386
rect 4072 11326 4098 11386
rect 3698 11324 3734 11326
rect 3798 11324 3822 11326
rect 3886 11324 3910 11326
rect 3974 11324 3998 11326
rect 4062 11324 4098 11326
rect 3698 11308 4098 11324
rect 10898 11388 11298 11404
rect 10898 11386 10934 11388
rect 10998 11386 11022 11388
rect 11086 11386 11110 11388
rect 11174 11386 11198 11388
rect 11262 11386 11298 11388
rect 10898 11326 10924 11386
rect 11272 11326 11298 11386
rect 10898 11324 10934 11326
rect 10998 11324 11022 11326
rect 11086 11324 11110 11326
rect 11174 11324 11198 11326
rect 11262 11324 11298 11326
rect 10898 11308 11298 11324
rect 18098 11388 18498 11404
rect 18098 11386 18134 11388
rect 18198 11386 18222 11388
rect 18286 11386 18310 11388
rect 18374 11386 18398 11388
rect 18462 11386 18498 11388
rect 18098 11326 18124 11386
rect 18472 11326 18498 11386
rect 18098 11324 18134 11326
rect 18198 11324 18222 11326
rect 18286 11324 18310 11326
rect 18374 11324 18398 11326
rect 18462 11324 18498 11326
rect 18098 11308 18498 11324
rect 25298 11388 25698 11404
rect 25298 11386 25334 11388
rect 25398 11386 25422 11388
rect 25486 11386 25510 11388
rect 25574 11386 25598 11388
rect 25662 11386 25698 11388
rect 25298 11326 25324 11386
rect 25672 11326 25698 11386
rect 25298 11324 25334 11326
rect 25398 11324 25422 11326
rect 25486 11324 25510 11326
rect 25574 11324 25598 11326
rect 25662 11324 25698 11326
rect 25298 11308 25698 11324
rect 32498 11387 32898 11404
rect 32498 11385 32534 11387
rect 32598 11385 32622 11387
rect 32686 11385 32710 11387
rect 32774 11385 32798 11387
rect 32862 11385 32898 11387
rect 32498 11325 32524 11385
rect 32872 11325 32898 11385
rect 32498 11323 32534 11325
rect 32598 11323 32622 11325
rect 32686 11323 32710 11325
rect 32774 11323 32798 11325
rect 32862 11323 32898 11325
rect 32498 11307 32898 11323
rect 36500 10748 36700 10908
rect 800 10332 1116 10470
rect 34364 9848 34680 9986
rect 3698 9212 4098 9228
rect 3698 9210 3734 9212
rect 3798 9210 3822 9212
rect 3886 9210 3910 9212
rect 3974 9210 3998 9212
rect 4062 9210 4098 9212
rect 3698 9150 3724 9210
rect 4072 9150 4098 9210
rect 3698 9148 3734 9150
rect 3798 9148 3822 9150
rect 3886 9148 3910 9150
rect 3974 9148 3998 9150
rect 4062 9148 4098 9150
rect 3698 9132 4098 9148
rect 10898 9212 11298 9228
rect 10898 9210 10934 9212
rect 10998 9210 11022 9212
rect 11086 9210 11110 9212
rect 11174 9210 11198 9212
rect 11262 9210 11298 9212
rect 10898 9150 10924 9210
rect 11272 9150 11298 9210
rect 10898 9148 10934 9150
rect 10998 9148 11022 9150
rect 11086 9148 11110 9150
rect 11174 9148 11198 9150
rect 11262 9148 11298 9150
rect 10898 9132 11298 9148
rect 18098 9212 18498 9228
rect 18098 9210 18134 9212
rect 18198 9210 18222 9212
rect 18286 9210 18310 9212
rect 18374 9210 18398 9212
rect 18462 9210 18498 9212
rect 18098 9150 18124 9210
rect 18472 9150 18498 9210
rect 18098 9148 18134 9150
rect 18198 9148 18222 9150
rect 18286 9148 18310 9150
rect 18374 9148 18398 9150
rect 18462 9148 18498 9150
rect 18098 9132 18498 9148
rect 25298 9212 25698 9228
rect 25298 9210 25334 9212
rect 25398 9210 25422 9212
rect 25486 9210 25510 9212
rect 25574 9210 25598 9212
rect 25662 9210 25698 9212
rect 25298 9150 25324 9210
rect 25672 9150 25698 9210
rect 25298 9148 25334 9150
rect 25398 9148 25422 9150
rect 25486 9148 25510 9150
rect 25574 9148 25598 9150
rect 25662 9148 25698 9150
rect 25298 9132 25698 9148
rect 32498 9212 32898 9228
rect 32498 9210 32534 9212
rect 32598 9210 32622 9212
rect 32686 9210 32710 9212
rect 32774 9210 32798 9212
rect 32862 9210 32898 9212
rect 32498 9150 32524 9210
rect 32872 9150 32898 9210
rect 32498 9148 32534 9150
rect 32598 9148 32622 9150
rect 32686 9148 32710 9150
rect 32774 9148 32798 9150
rect 32862 9148 32898 9150
rect 32498 9132 32898 9148
rect 3698 7036 4098 7052
rect 3698 7034 3734 7036
rect 3798 7034 3822 7036
rect 3886 7034 3910 7036
rect 3974 7034 3998 7036
rect 4062 7034 4098 7036
rect 3698 6974 3724 7034
rect 4072 6974 4098 7034
rect 3698 6972 3734 6974
rect 3798 6972 3822 6974
rect 3886 6972 3910 6974
rect 3974 6972 3998 6974
rect 4062 6972 4098 6974
rect 3698 6956 4098 6972
rect 10898 7036 11298 7052
rect 10898 7034 10934 7036
rect 10998 7034 11022 7036
rect 11086 7034 11110 7036
rect 11174 7034 11198 7036
rect 11262 7034 11298 7036
rect 10898 6974 10924 7034
rect 11272 6974 11298 7034
rect 10898 6972 10934 6974
rect 10998 6972 11022 6974
rect 11086 6972 11110 6974
rect 11174 6972 11198 6974
rect 11262 6972 11298 6974
rect 10898 6956 11298 6972
rect 25298 7036 25698 7052
rect 25298 7034 25334 7036
rect 25398 7034 25422 7036
rect 25486 7034 25510 7036
rect 25574 7034 25598 7036
rect 25662 7034 25698 7036
rect 25298 6974 25324 7034
rect 25672 6974 25698 7034
rect 25298 6972 25334 6974
rect 25398 6972 25422 6974
rect 25486 6972 25510 6974
rect 25574 6972 25598 6974
rect 25662 6972 25698 6974
rect 25298 6956 25698 6972
rect 32498 7036 32898 7052
rect 32498 7034 32534 7036
rect 32598 7034 32622 7036
rect 32686 7034 32710 7036
rect 32774 7034 32798 7036
rect 32862 7034 32898 7036
rect 32498 6974 32524 7034
rect 32872 6974 32898 7034
rect 32498 6972 32534 6974
rect 32598 6972 32622 6974
rect 32686 6972 32710 6974
rect 32774 6972 32798 6974
rect 32862 6972 32898 6974
rect 32498 6956 32898 6972
rect 2654 6202 2814 6402
rect 6254 6202 6414 6402
rect 12154 6202 12314 6402
rect 18054 6202 18214 6402
rect 23954 6202 24114 6402
rect 29854 6202 30014 6402
rect 33272 6202 33432 6402
rect 7298 6082 7698 6100
rect 7298 6080 7334 6082
rect 7398 6080 7422 6082
rect 7486 6080 7510 6082
rect 7574 6080 7598 6082
rect 7662 6080 7698 6082
rect 7298 6020 7324 6080
rect 7672 6020 7698 6080
rect 7298 6018 7334 6020
rect 7398 6018 7422 6020
rect 7486 6018 7510 6020
rect 7574 6018 7598 6020
rect 7662 6018 7698 6020
rect 7298 6000 7698 6018
rect 14498 6082 14898 6100
rect 14498 6080 14534 6082
rect 14598 6080 14622 6082
rect 14686 6080 14710 6082
rect 14774 6080 14798 6082
rect 14862 6080 14898 6082
rect 14498 6020 14524 6080
rect 14872 6020 14898 6080
rect 14498 6018 14534 6020
rect 14598 6018 14622 6020
rect 14686 6018 14710 6020
rect 14774 6018 14798 6020
rect 14862 6018 14898 6020
rect 14498 6000 14898 6018
rect 21698 6082 22098 6100
rect 21698 6080 21734 6082
rect 21798 6080 21822 6082
rect 21886 6080 21910 6082
rect 21974 6080 21998 6082
rect 22062 6080 22098 6082
rect 21698 6020 21724 6080
rect 22072 6020 22098 6080
rect 21698 6018 21734 6020
rect 21798 6018 21822 6020
rect 21886 6018 21910 6020
rect 21974 6018 21998 6020
rect 22062 6018 22098 6020
rect 21698 6000 22098 6018
rect 28898 6082 29298 6100
rect 28898 6080 28934 6082
rect 28998 6080 29022 6082
rect 29086 6080 29110 6082
rect 29174 6080 29198 6082
rect 29262 6080 29298 6082
rect 28898 6020 28924 6080
rect 29272 6020 29298 6080
rect 28898 6018 28934 6020
rect 28998 6018 29022 6020
rect 29086 6018 29110 6020
rect 29174 6018 29198 6020
rect 29262 6018 29298 6020
rect 28898 6000 29298 6018
<< via2 >>
rect 7334 14480 7398 14482
rect 7422 14480 7486 14482
rect 7510 14480 7574 14482
rect 7598 14480 7662 14482
rect 7334 14420 7384 14480
rect 7384 14420 7396 14480
rect 7396 14420 7398 14480
rect 7422 14420 7456 14480
rect 7456 14420 7468 14480
rect 7468 14420 7486 14480
rect 7510 14420 7528 14480
rect 7528 14420 7540 14480
rect 7540 14420 7574 14480
rect 7598 14420 7600 14480
rect 7600 14420 7612 14480
rect 7612 14420 7662 14480
rect 7334 14418 7398 14420
rect 7422 14418 7486 14420
rect 7510 14418 7574 14420
rect 7598 14418 7662 14420
rect 14534 14480 14598 14482
rect 14622 14480 14686 14482
rect 14710 14480 14774 14482
rect 14798 14480 14862 14482
rect 14534 14420 14584 14480
rect 14584 14420 14596 14480
rect 14596 14420 14598 14480
rect 14622 14420 14656 14480
rect 14656 14420 14668 14480
rect 14668 14420 14686 14480
rect 14710 14420 14728 14480
rect 14728 14420 14740 14480
rect 14740 14420 14774 14480
rect 14798 14420 14800 14480
rect 14800 14420 14812 14480
rect 14812 14420 14862 14480
rect 14534 14418 14598 14420
rect 14622 14418 14686 14420
rect 14710 14418 14774 14420
rect 14798 14418 14862 14420
rect 21734 14480 21798 14482
rect 21822 14480 21886 14482
rect 21910 14480 21974 14482
rect 21998 14480 22062 14482
rect 21734 14420 21784 14480
rect 21784 14420 21796 14480
rect 21796 14420 21798 14480
rect 21822 14420 21856 14480
rect 21856 14420 21868 14480
rect 21868 14420 21886 14480
rect 21910 14420 21928 14480
rect 21928 14420 21940 14480
rect 21940 14420 21974 14480
rect 21998 14420 22000 14480
rect 22000 14420 22012 14480
rect 22012 14420 22062 14480
rect 21734 14418 21798 14420
rect 21822 14418 21886 14420
rect 21910 14418 21974 14420
rect 21998 14418 22062 14420
rect 28934 14480 28998 14482
rect 29022 14480 29086 14482
rect 29110 14480 29174 14482
rect 29198 14480 29262 14482
rect 28934 14420 28984 14480
rect 28984 14420 28996 14480
rect 28996 14420 28998 14480
rect 29022 14420 29056 14480
rect 29056 14420 29068 14480
rect 29068 14420 29086 14480
rect 29110 14420 29128 14480
rect 29128 14420 29140 14480
rect 29140 14420 29174 14480
rect 29198 14420 29200 14480
rect 29200 14420 29212 14480
rect 29212 14420 29262 14480
rect 28934 14418 28998 14420
rect 29022 14418 29086 14420
rect 29110 14418 29174 14420
rect 29198 14418 29262 14420
rect 3734 13562 3798 13564
rect 3822 13562 3886 13564
rect 3910 13562 3974 13564
rect 3998 13562 4062 13564
rect 3734 13502 3784 13562
rect 3784 13502 3796 13562
rect 3796 13502 3798 13562
rect 3822 13502 3856 13562
rect 3856 13502 3868 13562
rect 3868 13502 3886 13562
rect 3910 13502 3928 13562
rect 3928 13502 3940 13562
rect 3940 13502 3974 13562
rect 3998 13502 4000 13562
rect 4000 13502 4012 13562
rect 4012 13502 4062 13562
rect 3734 13500 3798 13502
rect 3822 13500 3886 13502
rect 3910 13500 3974 13502
rect 3998 13500 4062 13502
rect 10934 13562 10998 13564
rect 11022 13562 11086 13564
rect 11110 13562 11174 13564
rect 11198 13562 11262 13564
rect 10934 13502 10984 13562
rect 10984 13502 10996 13562
rect 10996 13502 10998 13562
rect 11022 13502 11056 13562
rect 11056 13502 11068 13562
rect 11068 13502 11086 13562
rect 11110 13502 11128 13562
rect 11128 13502 11140 13562
rect 11140 13502 11174 13562
rect 11198 13502 11200 13562
rect 11200 13502 11212 13562
rect 11212 13502 11262 13562
rect 10934 13500 10998 13502
rect 11022 13500 11086 13502
rect 11110 13500 11174 13502
rect 11198 13500 11262 13502
rect 18134 13562 18198 13564
rect 18222 13562 18286 13564
rect 18310 13562 18374 13564
rect 18398 13562 18462 13564
rect 18134 13502 18184 13562
rect 18184 13502 18196 13562
rect 18196 13502 18198 13562
rect 18222 13502 18256 13562
rect 18256 13502 18268 13562
rect 18268 13502 18286 13562
rect 18310 13502 18328 13562
rect 18328 13502 18340 13562
rect 18340 13502 18374 13562
rect 18398 13502 18400 13562
rect 18400 13502 18412 13562
rect 18412 13502 18462 13562
rect 18134 13500 18198 13502
rect 18222 13500 18286 13502
rect 18310 13500 18374 13502
rect 18398 13500 18462 13502
rect 25334 13562 25398 13564
rect 25422 13562 25486 13564
rect 25510 13562 25574 13564
rect 25598 13562 25662 13564
rect 25334 13502 25384 13562
rect 25384 13502 25396 13562
rect 25396 13502 25398 13562
rect 25422 13502 25456 13562
rect 25456 13502 25468 13562
rect 25468 13502 25486 13562
rect 25510 13502 25528 13562
rect 25528 13502 25540 13562
rect 25540 13502 25574 13562
rect 25598 13502 25600 13562
rect 25600 13502 25612 13562
rect 25612 13502 25662 13562
rect 25334 13500 25398 13502
rect 25422 13500 25486 13502
rect 25510 13500 25574 13502
rect 25598 13500 25662 13502
rect 32534 13562 32598 13564
rect 32622 13562 32686 13564
rect 32710 13562 32774 13564
rect 32798 13562 32862 13564
rect 32534 13502 32584 13562
rect 32584 13502 32596 13562
rect 32596 13502 32598 13562
rect 32622 13502 32656 13562
rect 32656 13502 32668 13562
rect 32668 13502 32686 13562
rect 32710 13502 32728 13562
rect 32728 13502 32740 13562
rect 32740 13502 32774 13562
rect 32798 13502 32800 13562
rect 32800 13502 32812 13562
rect 32812 13502 32862 13562
rect 32534 13500 32598 13502
rect 32622 13500 32686 13502
rect 32710 13500 32774 13502
rect 32798 13500 32862 13502
rect 3734 12474 3798 12476
rect 3822 12474 3886 12476
rect 3910 12474 3974 12476
rect 3998 12474 4062 12476
rect 3734 12414 3784 12474
rect 3784 12414 3796 12474
rect 3796 12414 3798 12474
rect 3822 12414 3856 12474
rect 3856 12414 3868 12474
rect 3868 12414 3886 12474
rect 3910 12414 3928 12474
rect 3928 12414 3940 12474
rect 3940 12414 3974 12474
rect 3998 12414 4000 12474
rect 4000 12414 4012 12474
rect 4012 12414 4062 12474
rect 3734 12412 3798 12414
rect 3822 12412 3886 12414
rect 3910 12412 3974 12414
rect 3998 12412 4062 12414
rect 134 11930 198 11932
rect 222 11930 286 11932
rect 310 11930 374 11932
rect 398 11930 462 11932
rect 134 11870 184 11930
rect 184 11870 196 11930
rect 196 11870 198 11930
rect 222 11870 256 11930
rect 256 11870 268 11930
rect 268 11870 286 11930
rect 310 11870 328 11930
rect 328 11870 340 11930
rect 340 11870 374 11930
rect 398 11870 400 11930
rect 400 11870 412 11930
rect 412 11870 462 11930
rect 134 11868 198 11870
rect 222 11868 286 11870
rect 310 11868 374 11870
rect 398 11868 462 11870
rect 3734 11386 3798 11388
rect 3822 11386 3886 11388
rect 3910 11386 3974 11388
rect 3998 11386 4062 11388
rect 3734 11326 3784 11386
rect 3784 11326 3796 11386
rect 3796 11326 3798 11386
rect 3822 11326 3856 11386
rect 3856 11326 3868 11386
rect 3868 11326 3886 11386
rect 3910 11326 3928 11386
rect 3928 11326 3940 11386
rect 3940 11326 3974 11386
rect 3998 11326 4000 11386
rect 4000 11326 4012 11386
rect 4012 11326 4062 11386
rect 3734 11324 3798 11326
rect 3822 11324 3886 11326
rect 3910 11324 3974 11326
rect 3998 11324 4062 11326
rect 10934 11386 10998 11388
rect 11022 11386 11086 11388
rect 11110 11386 11174 11388
rect 11198 11386 11262 11388
rect 10934 11326 10984 11386
rect 10984 11326 10996 11386
rect 10996 11326 10998 11386
rect 11022 11326 11056 11386
rect 11056 11326 11068 11386
rect 11068 11326 11086 11386
rect 11110 11326 11128 11386
rect 11128 11326 11140 11386
rect 11140 11326 11174 11386
rect 11198 11326 11200 11386
rect 11200 11326 11212 11386
rect 11212 11326 11262 11386
rect 10934 11324 10998 11326
rect 11022 11324 11086 11326
rect 11110 11324 11174 11326
rect 11198 11324 11262 11326
rect 18134 11386 18198 11388
rect 18222 11386 18286 11388
rect 18310 11386 18374 11388
rect 18398 11386 18462 11388
rect 18134 11326 18184 11386
rect 18184 11326 18196 11386
rect 18196 11326 18198 11386
rect 18222 11326 18256 11386
rect 18256 11326 18268 11386
rect 18268 11326 18286 11386
rect 18310 11326 18328 11386
rect 18328 11326 18340 11386
rect 18340 11326 18374 11386
rect 18398 11326 18400 11386
rect 18400 11326 18412 11386
rect 18412 11326 18462 11386
rect 18134 11324 18198 11326
rect 18222 11324 18286 11326
rect 18310 11324 18374 11326
rect 18398 11324 18462 11326
rect 25334 11386 25398 11388
rect 25422 11386 25486 11388
rect 25510 11386 25574 11388
rect 25598 11386 25662 11388
rect 25334 11326 25384 11386
rect 25384 11326 25396 11386
rect 25396 11326 25398 11386
rect 25422 11326 25456 11386
rect 25456 11326 25468 11386
rect 25468 11326 25486 11386
rect 25510 11326 25528 11386
rect 25528 11326 25540 11386
rect 25540 11326 25574 11386
rect 25598 11326 25600 11386
rect 25600 11326 25612 11386
rect 25612 11326 25662 11386
rect 25334 11324 25398 11326
rect 25422 11324 25486 11326
rect 25510 11324 25574 11326
rect 25598 11324 25662 11326
rect 32534 11385 32598 11387
rect 32622 11385 32686 11387
rect 32710 11385 32774 11387
rect 32798 11385 32862 11387
rect 32534 11325 32584 11385
rect 32584 11325 32596 11385
rect 32596 11325 32598 11385
rect 32622 11325 32656 11385
rect 32656 11325 32668 11385
rect 32668 11325 32686 11385
rect 32710 11325 32728 11385
rect 32728 11325 32740 11385
rect 32740 11325 32774 11385
rect 32798 11325 32800 11385
rect 32800 11325 32812 11385
rect 32812 11325 32862 11385
rect 32534 11323 32598 11325
rect 32622 11323 32686 11325
rect 32710 11323 32774 11325
rect 32798 11323 32862 11325
rect 3734 9210 3798 9212
rect 3822 9210 3886 9212
rect 3910 9210 3974 9212
rect 3998 9210 4062 9212
rect 3734 9150 3784 9210
rect 3784 9150 3796 9210
rect 3796 9150 3798 9210
rect 3822 9150 3856 9210
rect 3856 9150 3868 9210
rect 3868 9150 3886 9210
rect 3910 9150 3928 9210
rect 3928 9150 3940 9210
rect 3940 9150 3974 9210
rect 3998 9150 4000 9210
rect 4000 9150 4012 9210
rect 4012 9150 4062 9210
rect 3734 9148 3798 9150
rect 3822 9148 3886 9150
rect 3910 9148 3974 9150
rect 3998 9148 4062 9150
rect 10934 9210 10998 9212
rect 11022 9210 11086 9212
rect 11110 9210 11174 9212
rect 11198 9210 11262 9212
rect 10934 9150 10984 9210
rect 10984 9150 10996 9210
rect 10996 9150 10998 9210
rect 11022 9150 11056 9210
rect 11056 9150 11068 9210
rect 11068 9150 11086 9210
rect 11110 9150 11128 9210
rect 11128 9150 11140 9210
rect 11140 9150 11174 9210
rect 11198 9150 11200 9210
rect 11200 9150 11212 9210
rect 11212 9150 11262 9210
rect 10934 9148 10998 9150
rect 11022 9148 11086 9150
rect 11110 9148 11174 9150
rect 11198 9148 11262 9150
rect 18134 9210 18198 9212
rect 18222 9210 18286 9212
rect 18310 9210 18374 9212
rect 18398 9210 18462 9212
rect 18134 9150 18184 9210
rect 18184 9150 18196 9210
rect 18196 9150 18198 9210
rect 18222 9150 18256 9210
rect 18256 9150 18268 9210
rect 18268 9150 18286 9210
rect 18310 9150 18328 9210
rect 18328 9150 18340 9210
rect 18340 9150 18374 9210
rect 18398 9150 18400 9210
rect 18400 9150 18412 9210
rect 18412 9150 18462 9210
rect 18134 9148 18198 9150
rect 18222 9148 18286 9150
rect 18310 9148 18374 9150
rect 18398 9148 18462 9150
rect 25334 9210 25398 9212
rect 25422 9210 25486 9212
rect 25510 9210 25574 9212
rect 25598 9210 25662 9212
rect 25334 9150 25384 9210
rect 25384 9150 25396 9210
rect 25396 9150 25398 9210
rect 25422 9150 25456 9210
rect 25456 9150 25468 9210
rect 25468 9150 25486 9210
rect 25510 9150 25528 9210
rect 25528 9150 25540 9210
rect 25540 9150 25574 9210
rect 25598 9150 25600 9210
rect 25600 9150 25612 9210
rect 25612 9150 25662 9210
rect 25334 9148 25398 9150
rect 25422 9148 25486 9150
rect 25510 9148 25574 9150
rect 25598 9148 25662 9150
rect 32534 9210 32598 9212
rect 32622 9210 32686 9212
rect 32710 9210 32774 9212
rect 32798 9210 32862 9212
rect 32534 9150 32584 9210
rect 32584 9150 32596 9210
rect 32596 9150 32598 9210
rect 32622 9150 32656 9210
rect 32656 9150 32668 9210
rect 32668 9150 32686 9210
rect 32710 9150 32728 9210
rect 32728 9150 32740 9210
rect 32740 9150 32774 9210
rect 32798 9150 32800 9210
rect 32800 9150 32812 9210
rect 32812 9150 32862 9210
rect 32534 9148 32598 9150
rect 32622 9148 32686 9150
rect 32710 9148 32774 9150
rect 32798 9148 32862 9150
rect 3734 7034 3798 7036
rect 3822 7034 3886 7036
rect 3910 7034 3974 7036
rect 3998 7034 4062 7036
rect 3734 6974 3784 7034
rect 3784 6974 3796 7034
rect 3796 6974 3798 7034
rect 3822 6974 3856 7034
rect 3856 6974 3868 7034
rect 3868 6974 3886 7034
rect 3910 6974 3928 7034
rect 3928 6974 3940 7034
rect 3940 6974 3974 7034
rect 3998 6974 4000 7034
rect 4000 6974 4012 7034
rect 4012 6974 4062 7034
rect 3734 6972 3798 6974
rect 3822 6972 3886 6974
rect 3910 6972 3974 6974
rect 3998 6972 4062 6974
rect 10934 7034 10998 7036
rect 11022 7034 11086 7036
rect 11110 7034 11174 7036
rect 11198 7034 11262 7036
rect 10934 6974 10984 7034
rect 10984 6974 10996 7034
rect 10996 6974 10998 7034
rect 11022 6974 11056 7034
rect 11056 6974 11068 7034
rect 11068 6974 11086 7034
rect 11110 6974 11128 7034
rect 11128 6974 11140 7034
rect 11140 6974 11174 7034
rect 11198 6974 11200 7034
rect 11200 6974 11212 7034
rect 11212 6974 11262 7034
rect 10934 6972 10998 6974
rect 11022 6972 11086 6974
rect 11110 6972 11174 6974
rect 11198 6972 11262 6974
rect 25334 7034 25398 7036
rect 25422 7034 25486 7036
rect 25510 7034 25574 7036
rect 25598 7034 25662 7036
rect 25334 6974 25384 7034
rect 25384 6974 25396 7034
rect 25396 6974 25398 7034
rect 25422 6974 25456 7034
rect 25456 6974 25468 7034
rect 25468 6974 25486 7034
rect 25510 6974 25528 7034
rect 25528 6974 25540 7034
rect 25540 6974 25574 7034
rect 25598 6974 25600 7034
rect 25600 6974 25612 7034
rect 25612 6974 25662 7034
rect 25334 6972 25398 6974
rect 25422 6972 25486 6974
rect 25510 6972 25574 6974
rect 25598 6972 25662 6974
rect 32534 7034 32598 7036
rect 32622 7034 32686 7036
rect 32710 7034 32774 7036
rect 32798 7034 32862 7036
rect 32534 6974 32584 7034
rect 32584 6974 32596 7034
rect 32596 6974 32598 7034
rect 32622 6974 32656 7034
rect 32656 6974 32668 7034
rect 32668 6974 32686 7034
rect 32710 6974 32728 7034
rect 32728 6974 32740 7034
rect 32740 6974 32774 7034
rect 32798 6974 32800 7034
rect 32800 6974 32812 7034
rect 32812 6974 32862 7034
rect 32534 6972 32598 6974
rect 32622 6972 32686 6974
rect 32710 6972 32774 6974
rect 32798 6972 32862 6974
rect 7334 6080 7398 6082
rect 7422 6080 7486 6082
rect 7510 6080 7574 6082
rect 7598 6080 7662 6082
rect 7334 6020 7384 6080
rect 7384 6020 7396 6080
rect 7396 6020 7398 6080
rect 7422 6020 7456 6080
rect 7456 6020 7468 6080
rect 7468 6020 7486 6080
rect 7510 6020 7528 6080
rect 7528 6020 7540 6080
rect 7540 6020 7574 6080
rect 7598 6020 7600 6080
rect 7600 6020 7612 6080
rect 7612 6020 7662 6080
rect 7334 6018 7398 6020
rect 7422 6018 7486 6020
rect 7510 6018 7574 6020
rect 7598 6018 7662 6020
rect 14534 6080 14598 6082
rect 14622 6080 14686 6082
rect 14710 6080 14774 6082
rect 14798 6080 14862 6082
rect 14534 6020 14584 6080
rect 14584 6020 14596 6080
rect 14596 6020 14598 6080
rect 14622 6020 14656 6080
rect 14656 6020 14668 6080
rect 14668 6020 14686 6080
rect 14710 6020 14728 6080
rect 14728 6020 14740 6080
rect 14740 6020 14774 6080
rect 14798 6020 14800 6080
rect 14800 6020 14812 6080
rect 14812 6020 14862 6080
rect 14534 6018 14598 6020
rect 14622 6018 14686 6020
rect 14710 6018 14774 6020
rect 14798 6018 14862 6020
rect 21734 6080 21798 6082
rect 21822 6080 21886 6082
rect 21910 6080 21974 6082
rect 21998 6080 22062 6082
rect 21734 6020 21784 6080
rect 21784 6020 21796 6080
rect 21796 6020 21798 6080
rect 21822 6020 21856 6080
rect 21856 6020 21868 6080
rect 21868 6020 21886 6080
rect 21910 6020 21928 6080
rect 21928 6020 21940 6080
rect 21940 6020 21974 6080
rect 21998 6020 22000 6080
rect 22000 6020 22012 6080
rect 22012 6020 22062 6080
rect 21734 6018 21798 6020
rect 21822 6018 21886 6020
rect 21910 6018 21974 6020
rect 21998 6018 22062 6020
rect 28934 6080 28998 6082
rect 29022 6080 29086 6082
rect 29110 6080 29174 6082
rect 29198 6080 29262 6082
rect 28934 6020 28984 6080
rect 28984 6020 28996 6080
rect 28996 6020 28998 6080
rect 29022 6020 29056 6080
rect 29056 6020 29068 6080
rect 29068 6020 29086 6080
rect 29110 6020 29128 6080
rect 29128 6020 29140 6080
rect 29140 6020 29174 6080
rect 29198 6020 29200 6080
rect 29200 6020 29212 6080
rect 29212 6020 29262 6080
rect 28934 6018 28998 6020
rect 29022 6018 29086 6020
rect 29110 6018 29174 6020
rect 29198 6018 29262 6020
<< metal3 >>
rect 30800 21800 31800 22200
rect 30800 20600 31800 21000
rect 7298 14487 7698 14500
rect 7298 14414 7330 14487
rect 7402 14414 7418 14487
rect 7490 14414 7506 14487
rect 7578 14414 7594 14487
rect 7666 14414 7698 14487
rect 7298 14400 7698 14414
rect 14498 14487 14898 14500
rect 14498 14414 14530 14487
rect 14602 14414 14618 14487
rect 14690 14414 14706 14487
rect 14778 14414 14794 14487
rect 14866 14414 14898 14487
rect 14498 14400 14898 14414
rect 21698 14487 22098 14500
rect 21698 14414 21730 14487
rect 21802 14414 21818 14487
rect 21890 14414 21906 14487
rect 21978 14414 21994 14487
rect 22066 14414 22098 14487
rect 21698 14400 22098 14414
rect 28898 14487 29298 14500
rect 28898 14414 28930 14487
rect 29002 14414 29018 14487
rect 29090 14414 29106 14487
rect 29178 14414 29194 14487
rect 29266 14414 29298 14487
rect 28898 14400 29298 14414
rect 3698 13568 4098 13580
rect 3698 13496 3730 13568
rect 3802 13496 3818 13568
rect 3890 13496 3906 13568
rect 3978 13496 3994 13568
rect 4066 13496 4098 13568
rect 3698 13484 4098 13496
rect 10898 13568 11298 13580
rect 10898 13496 10930 13568
rect 11002 13496 11018 13568
rect 11090 13496 11106 13568
rect 11178 13496 11194 13568
rect 11266 13496 11298 13568
rect 10898 13484 11298 13496
rect 18098 13568 18498 13580
rect 18098 13496 18130 13568
rect 18202 13496 18218 13568
rect 18290 13496 18306 13568
rect 18378 13496 18394 13568
rect 18466 13496 18498 13568
rect 18098 13484 18498 13496
rect 25298 13568 25698 13580
rect 25298 13496 25330 13568
rect 25402 13496 25418 13568
rect 25490 13496 25506 13568
rect 25578 13496 25594 13568
rect 25666 13496 25698 13568
rect 25298 13484 25698 13496
rect 32498 13568 32898 13580
rect 32498 13496 32530 13568
rect 32602 13496 32618 13568
rect 32690 13496 32706 13568
rect 32778 13496 32794 13568
rect 32866 13496 32898 13568
rect 32498 13484 32898 13496
rect 3698 12480 4098 12492
rect 3698 12408 3730 12480
rect 3802 12408 3818 12480
rect 3890 12408 3906 12480
rect 3978 12408 3994 12480
rect 4066 12408 4098 12480
rect 3698 12396 4098 12408
rect 98 11937 498 11948
rect 98 11864 130 11937
rect 202 11864 218 11937
rect 290 11864 306 11937
rect 378 11864 394 11937
rect 466 11864 498 11937
rect 98 11852 498 11864
rect 3698 11392 4098 11404
rect 3698 11320 3730 11392
rect 3802 11320 3818 11392
rect 3890 11320 3906 11392
rect 3978 11320 3994 11392
rect 4066 11320 4098 11392
rect 3698 11308 4098 11320
rect 10898 11392 11298 11404
rect 10898 11320 10930 11392
rect 11002 11320 11018 11392
rect 11090 11320 11106 11392
rect 11178 11320 11194 11392
rect 11266 11320 11298 11392
rect 10898 11308 11298 11320
rect 18098 11392 18498 11404
rect 18098 11320 18130 11392
rect 18202 11320 18218 11392
rect 18290 11320 18306 11392
rect 18378 11320 18394 11392
rect 18466 11320 18498 11392
rect 18098 11308 18498 11320
rect 25298 11392 25698 11404
rect 25298 11320 25330 11392
rect 25402 11320 25418 11392
rect 25490 11320 25506 11392
rect 25578 11320 25594 11392
rect 25666 11320 25698 11392
rect 25298 11308 25698 11320
rect 32498 11392 32898 11404
rect 32498 11319 32530 11392
rect 32602 11319 32618 11392
rect 32690 11319 32706 11392
rect 32778 11319 32794 11392
rect 32866 11319 32898 11392
rect 32498 11307 32898 11319
rect 3698 9217 4098 9228
rect 3698 9144 3730 9217
rect 3802 9144 3818 9217
rect 3890 9144 3906 9217
rect 3978 9144 3994 9217
rect 4066 9144 4098 9217
rect 3698 9132 4098 9144
rect 10898 9217 11298 9228
rect 10898 9144 10930 9217
rect 11002 9144 11018 9217
rect 11090 9144 11106 9217
rect 11178 9144 11194 9217
rect 11266 9144 11298 9217
rect 10898 9132 11298 9144
rect 18098 9217 18498 9228
rect 18098 9144 18130 9217
rect 18202 9144 18218 9217
rect 18290 9144 18306 9217
rect 18378 9144 18394 9217
rect 18466 9144 18498 9217
rect 18098 9132 18498 9144
rect 25298 9217 25698 9228
rect 25298 9144 25330 9217
rect 25402 9144 25418 9217
rect 25490 9144 25506 9217
rect 25578 9144 25594 9217
rect 25666 9144 25698 9217
rect 25298 9132 25698 9144
rect 32498 9217 32898 9228
rect 32498 9144 32530 9217
rect 32602 9144 32618 9217
rect 32690 9144 32706 9217
rect 32778 9144 32794 9217
rect 32866 9144 32898 9217
rect 32498 9132 32898 9144
rect 3698 7041 4098 7052
rect 3698 6968 3730 7041
rect 3802 6968 3818 7041
rect 3890 6968 3906 7041
rect 3978 6968 3994 7041
rect 4066 6968 4098 7041
rect 3698 6956 4098 6968
rect 10898 7041 11298 7052
rect 10898 6968 10930 7041
rect 11002 6968 11018 7041
rect 11090 6968 11106 7041
rect 11178 6968 11194 7041
rect 11266 6968 11298 7041
rect 10898 6956 11298 6968
rect 25298 7041 25698 7052
rect 25298 6968 25330 7041
rect 25402 6968 25418 7041
rect 25490 6968 25506 7041
rect 25578 6968 25594 7041
rect 25666 6968 25698 7041
rect 25298 6956 25698 6968
rect 32498 7041 32898 7052
rect 32498 6968 32530 7041
rect 32602 6968 32618 7041
rect 32690 6968 32706 7041
rect 32778 6968 32794 7041
rect 32866 6968 32898 7041
rect 32498 6956 32898 6968
rect 7298 6087 7698 6100
rect 7298 6014 7330 6087
rect 7402 6014 7418 6087
rect 7490 6014 7506 6087
rect 7578 6014 7594 6087
rect 7666 6014 7698 6087
rect 7298 6000 7698 6014
rect 14498 6087 14898 6100
rect 14498 6014 14530 6087
rect 14602 6014 14618 6087
rect 14690 6014 14706 6087
rect 14778 6014 14794 6087
rect 14866 6014 14898 6087
rect 14498 6000 14898 6014
rect 21698 6087 22098 6100
rect 21698 6014 21730 6087
rect 21802 6014 21818 6087
rect 21890 6014 21906 6087
rect 21978 6014 21994 6087
rect 22066 6014 22098 6087
rect 21698 6000 22098 6014
rect 28898 6087 29298 6100
rect 28898 6014 28930 6087
rect 29002 6014 29018 6087
rect 29090 6014 29106 6087
rect 29178 6014 29194 6087
rect 29266 6014 29298 6087
rect 28898 6000 29298 6014
<< via3 >>
rect 7330 14482 7402 14487
rect 7330 14418 7334 14482
rect 7334 14418 7398 14482
rect 7398 14418 7402 14482
rect 7330 14414 7402 14418
rect 7418 14482 7490 14487
rect 7418 14418 7422 14482
rect 7422 14418 7486 14482
rect 7486 14418 7490 14482
rect 7418 14414 7490 14418
rect 7506 14482 7578 14487
rect 7506 14418 7510 14482
rect 7510 14418 7574 14482
rect 7574 14418 7578 14482
rect 7506 14414 7578 14418
rect 7594 14482 7666 14487
rect 7594 14418 7598 14482
rect 7598 14418 7662 14482
rect 7662 14418 7666 14482
rect 7594 14414 7666 14418
rect 14530 14482 14602 14487
rect 14530 14418 14534 14482
rect 14534 14418 14598 14482
rect 14598 14418 14602 14482
rect 14530 14414 14602 14418
rect 14618 14482 14690 14487
rect 14618 14418 14622 14482
rect 14622 14418 14686 14482
rect 14686 14418 14690 14482
rect 14618 14414 14690 14418
rect 14706 14482 14778 14487
rect 14706 14418 14710 14482
rect 14710 14418 14774 14482
rect 14774 14418 14778 14482
rect 14706 14414 14778 14418
rect 14794 14482 14866 14487
rect 14794 14418 14798 14482
rect 14798 14418 14862 14482
rect 14862 14418 14866 14482
rect 14794 14414 14866 14418
rect 21730 14482 21802 14487
rect 21730 14418 21734 14482
rect 21734 14418 21798 14482
rect 21798 14418 21802 14482
rect 21730 14414 21802 14418
rect 21818 14482 21890 14487
rect 21818 14418 21822 14482
rect 21822 14418 21886 14482
rect 21886 14418 21890 14482
rect 21818 14414 21890 14418
rect 21906 14482 21978 14487
rect 21906 14418 21910 14482
rect 21910 14418 21974 14482
rect 21974 14418 21978 14482
rect 21906 14414 21978 14418
rect 21994 14482 22066 14487
rect 21994 14418 21998 14482
rect 21998 14418 22062 14482
rect 22062 14418 22066 14482
rect 21994 14414 22066 14418
rect 28930 14482 29002 14487
rect 28930 14418 28934 14482
rect 28934 14418 28998 14482
rect 28998 14418 29002 14482
rect 28930 14414 29002 14418
rect 29018 14482 29090 14487
rect 29018 14418 29022 14482
rect 29022 14418 29086 14482
rect 29086 14418 29090 14482
rect 29018 14414 29090 14418
rect 29106 14482 29178 14487
rect 29106 14418 29110 14482
rect 29110 14418 29174 14482
rect 29174 14418 29178 14482
rect 29106 14414 29178 14418
rect 29194 14482 29266 14487
rect 29194 14418 29198 14482
rect 29198 14418 29262 14482
rect 29262 14418 29266 14482
rect 29194 14414 29266 14418
rect 3730 13564 3802 13568
rect 3730 13500 3734 13564
rect 3734 13500 3798 13564
rect 3798 13500 3802 13564
rect 3730 13496 3802 13500
rect 3818 13564 3890 13568
rect 3818 13500 3822 13564
rect 3822 13500 3886 13564
rect 3886 13500 3890 13564
rect 3818 13496 3890 13500
rect 3906 13564 3978 13568
rect 3906 13500 3910 13564
rect 3910 13500 3974 13564
rect 3974 13500 3978 13564
rect 3906 13496 3978 13500
rect 3994 13564 4066 13568
rect 3994 13500 3998 13564
rect 3998 13500 4062 13564
rect 4062 13500 4066 13564
rect 3994 13496 4066 13500
rect 10930 13564 11002 13568
rect 10930 13500 10934 13564
rect 10934 13500 10998 13564
rect 10998 13500 11002 13564
rect 10930 13496 11002 13500
rect 11018 13564 11090 13568
rect 11018 13500 11022 13564
rect 11022 13500 11086 13564
rect 11086 13500 11090 13564
rect 11018 13496 11090 13500
rect 11106 13564 11178 13568
rect 11106 13500 11110 13564
rect 11110 13500 11174 13564
rect 11174 13500 11178 13564
rect 11106 13496 11178 13500
rect 11194 13564 11266 13568
rect 11194 13500 11198 13564
rect 11198 13500 11262 13564
rect 11262 13500 11266 13564
rect 11194 13496 11266 13500
rect 18130 13564 18202 13568
rect 18130 13500 18134 13564
rect 18134 13500 18198 13564
rect 18198 13500 18202 13564
rect 18130 13496 18202 13500
rect 18218 13564 18290 13568
rect 18218 13500 18222 13564
rect 18222 13500 18286 13564
rect 18286 13500 18290 13564
rect 18218 13496 18290 13500
rect 18306 13564 18378 13568
rect 18306 13500 18310 13564
rect 18310 13500 18374 13564
rect 18374 13500 18378 13564
rect 18306 13496 18378 13500
rect 18394 13564 18466 13568
rect 18394 13500 18398 13564
rect 18398 13500 18462 13564
rect 18462 13500 18466 13564
rect 18394 13496 18466 13500
rect 25330 13564 25402 13568
rect 25330 13500 25334 13564
rect 25334 13500 25398 13564
rect 25398 13500 25402 13564
rect 25330 13496 25402 13500
rect 25418 13564 25490 13568
rect 25418 13500 25422 13564
rect 25422 13500 25486 13564
rect 25486 13500 25490 13564
rect 25418 13496 25490 13500
rect 25506 13564 25578 13568
rect 25506 13500 25510 13564
rect 25510 13500 25574 13564
rect 25574 13500 25578 13564
rect 25506 13496 25578 13500
rect 25594 13564 25666 13568
rect 25594 13500 25598 13564
rect 25598 13500 25662 13564
rect 25662 13500 25666 13564
rect 25594 13496 25666 13500
rect 32530 13564 32602 13568
rect 32530 13500 32534 13564
rect 32534 13500 32598 13564
rect 32598 13500 32602 13564
rect 32530 13496 32602 13500
rect 32618 13564 32690 13568
rect 32618 13500 32622 13564
rect 32622 13500 32686 13564
rect 32686 13500 32690 13564
rect 32618 13496 32690 13500
rect 32706 13564 32778 13568
rect 32706 13500 32710 13564
rect 32710 13500 32774 13564
rect 32774 13500 32778 13564
rect 32706 13496 32778 13500
rect 32794 13564 32866 13568
rect 32794 13500 32798 13564
rect 32798 13500 32862 13564
rect 32862 13500 32866 13564
rect 32794 13496 32866 13500
rect 3730 12476 3802 12480
rect 3730 12412 3734 12476
rect 3734 12412 3798 12476
rect 3798 12412 3802 12476
rect 3730 12408 3802 12412
rect 3818 12476 3890 12480
rect 3818 12412 3822 12476
rect 3822 12412 3886 12476
rect 3886 12412 3890 12476
rect 3818 12408 3890 12412
rect 3906 12476 3978 12480
rect 3906 12412 3910 12476
rect 3910 12412 3974 12476
rect 3974 12412 3978 12476
rect 3906 12408 3978 12412
rect 3994 12476 4066 12480
rect 3994 12412 3998 12476
rect 3998 12412 4062 12476
rect 4062 12412 4066 12476
rect 3994 12408 4066 12412
rect 130 11932 202 11937
rect 130 11868 134 11932
rect 134 11868 198 11932
rect 198 11868 202 11932
rect 130 11864 202 11868
rect 218 11932 290 11937
rect 218 11868 222 11932
rect 222 11868 286 11932
rect 286 11868 290 11932
rect 218 11864 290 11868
rect 306 11932 378 11937
rect 306 11868 310 11932
rect 310 11868 374 11932
rect 374 11868 378 11932
rect 306 11864 378 11868
rect 394 11932 466 11937
rect 394 11868 398 11932
rect 398 11868 462 11932
rect 462 11868 466 11932
rect 394 11864 466 11868
rect 3730 11388 3802 11392
rect 3730 11324 3734 11388
rect 3734 11324 3798 11388
rect 3798 11324 3802 11388
rect 3730 11320 3802 11324
rect 3818 11388 3890 11392
rect 3818 11324 3822 11388
rect 3822 11324 3886 11388
rect 3886 11324 3890 11388
rect 3818 11320 3890 11324
rect 3906 11388 3978 11392
rect 3906 11324 3910 11388
rect 3910 11324 3974 11388
rect 3974 11324 3978 11388
rect 3906 11320 3978 11324
rect 3994 11388 4066 11392
rect 3994 11324 3998 11388
rect 3998 11324 4062 11388
rect 4062 11324 4066 11388
rect 3994 11320 4066 11324
rect 10930 11388 11002 11392
rect 10930 11324 10934 11388
rect 10934 11324 10998 11388
rect 10998 11324 11002 11388
rect 10930 11320 11002 11324
rect 11018 11388 11090 11392
rect 11018 11324 11022 11388
rect 11022 11324 11086 11388
rect 11086 11324 11090 11388
rect 11018 11320 11090 11324
rect 11106 11388 11178 11392
rect 11106 11324 11110 11388
rect 11110 11324 11174 11388
rect 11174 11324 11178 11388
rect 11106 11320 11178 11324
rect 11194 11388 11266 11392
rect 11194 11324 11198 11388
rect 11198 11324 11262 11388
rect 11262 11324 11266 11388
rect 11194 11320 11266 11324
rect 18130 11388 18202 11392
rect 18130 11324 18134 11388
rect 18134 11324 18198 11388
rect 18198 11324 18202 11388
rect 18130 11320 18202 11324
rect 18218 11388 18290 11392
rect 18218 11324 18222 11388
rect 18222 11324 18286 11388
rect 18286 11324 18290 11388
rect 18218 11320 18290 11324
rect 18306 11388 18378 11392
rect 18306 11324 18310 11388
rect 18310 11324 18374 11388
rect 18374 11324 18378 11388
rect 18306 11320 18378 11324
rect 18394 11388 18466 11392
rect 18394 11324 18398 11388
rect 18398 11324 18462 11388
rect 18462 11324 18466 11388
rect 18394 11320 18466 11324
rect 25330 11388 25402 11392
rect 25330 11324 25334 11388
rect 25334 11324 25398 11388
rect 25398 11324 25402 11388
rect 25330 11320 25402 11324
rect 25418 11388 25490 11392
rect 25418 11324 25422 11388
rect 25422 11324 25486 11388
rect 25486 11324 25490 11388
rect 25418 11320 25490 11324
rect 25506 11388 25578 11392
rect 25506 11324 25510 11388
rect 25510 11324 25574 11388
rect 25574 11324 25578 11388
rect 25506 11320 25578 11324
rect 25594 11388 25666 11392
rect 25594 11324 25598 11388
rect 25598 11324 25662 11388
rect 25662 11324 25666 11388
rect 25594 11320 25666 11324
rect 32530 11387 32602 11392
rect 32530 11323 32534 11387
rect 32534 11323 32598 11387
rect 32598 11323 32602 11387
rect 32530 11319 32602 11323
rect 32618 11387 32690 11392
rect 32618 11323 32622 11387
rect 32622 11323 32686 11387
rect 32686 11323 32690 11387
rect 32618 11319 32690 11323
rect 32706 11387 32778 11392
rect 32706 11323 32710 11387
rect 32710 11323 32774 11387
rect 32774 11323 32778 11387
rect 32706 11319 32778 11323
rect 32794 11387 32866 11392
rect 32794 11323 32798 11387
rect 32798 11323 32862 11387
rect 32862 11323 32866 11387
rect 32794 11319 32866 11323
rect 3730 9212 3802 9217
rect 3730 9148 3734 9212
rect 3734 9148 3798 9212
rect 3798 9148 3802 9212
rect 3730 9144 3802 9148
rect 3818 9212 3890 9217
rect 3818 9148 3822 9212
rect 3822 9148 3886 9212
rect 3886 9148 3890 9212
rect 3818 9144 3890 9148
rect 3906 9212 3978 9217
rect 3906 9148 3910 9212
rect 3910 9148 3974 9212
rect 3974 9148 3978 9212
rect 3906 9144 3978 9148
rect 3994 9212 4066 9217
rect 3994 9148 3998 9212
rect 3998 9148 4062 9212
rect 4062 9148 4066 9212
rect 3994 9144 4066 9148
rect 10930 9212 11002 9217
rect 10930 9148 10934 9212
rect 10934 9148 10998 9212
rect 10998 9148 11002 9212
rect 10930 9144 11002 9148
rect 11018 9212 11090 9217
rect 11018 9148 11022 9212
rect 11022 9148 11086 9212
rect 11086 9148 11090 9212
rect 11018 9144 11090 9148
rect 11106 9212 11178 9217
rect 11106 9148 11110 9212
rect 11110 9148 11174 9212
rect 11174 9148 11178 9212
rect 11106 9144 11178 9148
rect 11194 9212 11266 9217
rect 11194 9148 11198 9212
rect 11198 9148 11262 9212
rect 11262 9148 11266 9212
rect 11194 9144 11266 9148
rect 18130 9212 18202 9217
rect 18130 9148 18134 9212
rect 18134 9148 18198 9212
rect 18198 9148 18202 9212
rect 18130 9144 18202 9148
rect 18218 9212 18290 9217
rect 18218 9148 18222 9212
rect 18222 9148 18286 9212
rect 18286 9148 18290 9212
rect 18218 9144 18290 9148
rect 18306 9212 18378 9217
rect 18306 9148 18310 9212
rect 18310 9148 18374 9212
rect 18374 9148 18378 9212
rect 18306 9144 18378 9148
rect 18394 9212 18466 9217
rect 18394 9148 18398 9212
rect 18398 9148 18462 9212
rect 18462 9148 18466 9212
rect 18394 9144 18466 9148
rect 25330 9212 25402 9217
rect 25330 9148 25334 9212
rect 25334 9148 25398 9212
rect 25398 9148 25402 9212
rect 25330 9144 25402 9148
rect 25418 9212 25490 9217
rect 25418 9148 25422 9212
rect 25422 9148 25486 9212
rect 25486 9148 25490 9212
rect 25418 9144 25490 9148
rect 25506 9212 25578 9217
rect 25506 9148 25510 9212
rect 25510 9148 25574 9212
rect 25574 9148 25578 9212
rect 25506 9144 25578 9148
rect 25594 9212 25666 9217
rect 25594 9148 25598 9212
rect 25598 9148 25662 9212
rect 25662 9148 25666 9212
rect 25594 9144 25666 9148
rect 32530 9212 32602 9217
rect 32530 9148 32534 9212
rect 32534 9148 32598 9212
rect 32598 9148 32602 9212
rect 32530 9144 32602 9148
rect 32618 9212 32690 9217
rect 32618 9148 32622 9212
rect 32622 9148 32686 9212
rect 32686 9148 32690 9212
rect 32618 9144 32690 9148
rect 32706 9212 32778 9217
rect 32706 9148 32710 9212
rect 32710 9148 32774 9212
rect 32774 9148 32778 9212
rect 32706 9144 32778 9148
rect 32794 9212 32866 9217
rect 32794 9148 32798 9212
rect 32798 9148 32862 9212
rect 32862 9148 32866 9212
rect 32794 9144 32866 9148
rect 3730 7036 3802 7041
rect 3730 6972 3734 7036
rect 3734 6972 3798 7036
rect 3798 6972 3802 7036
rect 3730 6968 3802 6972
rect 3818 7036 3890 7041
rect 3818 6972 3822 7036
rect 3822 6972 3886 7036
rect 3886 6972 3890 7036
rect 3818 6968 3890 6972
rect 3906 7036 3978 7041
rect 3906 6972 3910 7036
rect 3910 6972 3974 7036
rect 3974 6972 3978 7036
rect 3906 6968 3978 6972
rect 3994 7036 4066 7041
rect 3994 6972 3998 7036
rect 3998 6972 4062 7036
rect 4062 6972 4066 7036
rect 3994 6968 4066 6972
rect 10930 7036 11002 7041
rect 10930 6972 10934 7036
rect 10934 6972 10998 7036
rect 10998 6972 11002 7036
rect 10930 6968 11002 6972
rect 11018 7036 11090 7041
rect 11018 6972 11022 7036
rect 11022 6972 11086 7036
rect 11086 6972 11090 7036
rect 11018 6968 11090 6972
rect 11106 7036 11178 7041
rect 11106 6972 11110 7036
rect 11110 6972 11174 7036
rect 11174 6972 11178 7036
rect 11106 6968 11178 6972
rect 11194 7036 11266 7041
rect 11194 6972 11198 7036
rect 11198 6972 11262 7036
rect 11262 6972 11266 7036
rect 11194 6968 11266 6972
rect 25330 7036 25402 7041
rect 25330 6972 25334 7036
rect 25334 6972 25398 7036
rect 25398 6972 25402 7036
rect 25330 6968 25402 6972
rect 25418 7036 25490 7041
rect 25418 6972 25422 7036
rect 25422 6972 25486 7036
rect 25486 6972 25490 7036
rect 25418 6968 25490 6972
rect 25506 7036 25578 7041
rect 25506 6972 25510 7036
rect 25510 6972 25574 7036
rect 25574 6972 25578 7036
rect 25506 6968 25578 6972
rect 25594 7036 25666 7041
rect 25594 6972 25598 7036
rect 25598 6972 25662 7036
rect 25662 6972 25666 7036
rect 25594 6968 25666 6972
rect 32530 7036 32602 7041
rect 32530 6972 32534 7036
rect 32534 6972 32598 7036
rect 32598 6972 32602 7036
rect 32530 6968 32602 6972
rect 32618 7036 32690 7041
rect 32618 6972 32622 7036
rect 32622 6972 32686 7036
rect 32686 6972 32690 7036
rect 32618 6968 32690 6972
rect 32706 7036 32778 7041
rect 32706 6972 32710 7036
rect 32710 6972 32774 7036
rect 32774 6972 32778 7036
rect 32706 6968 32778 6972
rect 32794 7036 32866 7041
rect 32794 6972 32798 7036
rect 32798 6972 32862 7036
rect 32862 6972 32866 7036
rect 32794 6968 32866 6972
rect 7330 6082 7402 6087
rect 7330 6018 7334 6082
rect 7334 6018 7398 6082
rect 7398 6018 7402 6082
rect 7330 6014 7402 6018
rect 7418 6082 7490 6087
rect 7418 6018 7422 6082
rect 7422 6018 7486 6082
rect 7486 6018 7490 6082
rect 7418 6014 7490 6018
rect 7506 6082 7578 6087
rect 7506 6018 7510 6082
rect 7510 6018 7574 6082
rect 7574 6018 7578 6082
rect 7506 6014 7578 6018
rect 7594 6082 7666 6087
rect 7594 6018 7598 6082
rect 7598 6018 7662 6082
rect 7662 6018 7666 6082
rect 7594 6014 7666 6018
rect 14530 6082 14602 6087
rect 14530 6018 14534 6082
rect 14534 6018 14598 6082
rect 14598 6018 14602 6082
rect 14530 6014 14602 6018
rect 14618 6082 14690 6087
rect 14618 6018 14622 6082
rect 14622 6018 14686 6082
rect 14686 6018 14690 6082
rect 14618 6014 14690 6018
rect 14706 6082 14778 6087
rect 14706 6018 14710 6082
rect 14710 6018 14774 6082
rect 14774 6018 14778 6082
rect 14706 6014 14778 6018
rect 14794 6082 14866 6087
rect 14794 6018 14798 6082
rect 14798 6018 14862 6082
rect 14862 6018 14866 6082
rect 14794 6014 14866 6018
rect 21730 6082 21802 6087
rect 21730 6018 21734 6082
rect 21734 6018 21798 6082
rect 21798 6018 21802 6082
rect 21730 6014 21802 6018
rect 21818 6082 21890 6087
rect 21818 6018 21822 6082
rect 21822 6018 21886 6082
rect 21886 6018 21890 6082
rect 21818 6014 21890 6018
rect 21906 6082 21978 6087
rect 21906 6018 21910 6082
rect 21910 6018 21974 6082
rect 21974 6018 21978 6082
rect 21906 6014 21978 6018
rect 21994 6082 22066 6087
rect 21994 6018 21998 6082
rect 21998 6018 22062 6082
rect 22062 6018 22066 6082
rect 21994 6014 22066 6018
rect 28930 6082 29002 6087
rect 28930 6018 28934 6082
rect 28934 6018 28998 6082
rect 28998 6018 29002 6082
rect 28930 6014 29002 6018
rect 29018 6082 29090 6087
rect 29018 6018 29022 6082
rect 29022 6018 29086 6082
rect 29086 6018 29090 6082
rect 29018 6014 29090 6018
rect 29106 6082 29178 6087
rect 29106 6018 29110 6082
rect 29110 6018 29174 6082
rect 29174 6018 29178 6082
rect 29106 6014 29178 6018
rect 29194 6082 29266 6087
rect 29194 6018 29198 6082
rect 29198 6018 29262 6082
rect 29262 6018 29266 6082
rect 29194 6014 29266 6018
<< metal4 >>
rect 7298 14487 7698 14500
rect 7298 14414 7330 14487
rect 7402 14414 7418 14487
rect 7490 14414 7506 14487
rect 7578 14414 7594 14487
rect 7666 14414 7698 14487
rect 7298 14400 7698 14414
rect 14498 14487 14898 14500
rect 14498 14414 14530 14487
rect 14602 14414 14618 14487
rect 14690 14414 14706 14487
rect 14778 14414 14794 14487
rect 14866 14414 14898 14487
rect 14498 14400 14898 14414
rect 21698 14487 22098 14500
rect 21698 14414 21730 14487
rect 21802 14414 21818 14487
rect 21890 14414 21906 14487
rect 21978 14414 21994 14487
rect 22066 14414 22098 14487
rect 21698 14400 22098 14414
rect 28898 14487 29298 14500
rect 28898 14414 28930 14487
rect 29002 14414 29018 14487
rect 29090 14414 29106 14487
rect 29178 14414 29194 14487
rect 29266 14414 29298 14487
rect 28898 14400 29298 14414
rect 3698 13568 4098 13580
rect 3698 13496 3730 13568
rect 3802 13496 3818 13568
rect 3890 13496 3906 13568
rect 3978 13496 3994 13568
rect 4066 13496 4098 13568
rect 3698 13484 4098 13496
rect 10898 13568 11298 13580
rect 10898 13496 10930 13568
rect 11002 13496 11018 13568
rect 11090 13496 11106 13568
rect 11178 13496 11194 13568
rect 11266 13496 11298 13568
rect 10898 13484 11298 13496
rect 18098 13568 18498 13580
rect 18098 13496 18130 13568
rect 18202 13496 18218 13568
rect 18290 13496 18306 13568
rect 18378 13496 18394 13568
rect 18466 13496 18498 13568
rect 18098 13484 18498 13496
rect 25298 13568 25698 13580
rect 25298 13496 25330 13568
rect 25402 13496 25418 13568
rect 25490 13496 25506 13568
rect 25578 13496 25594 13568
rect 25666 13496 25698 13568
rect 25298 13484 25698 13496
rect 32498 13568 32898 13580
rect 32498 13496 32530 13568
rect 32602 13496 32618 13568
rect 32690 13496 32706 13568
rect 32778 13496 32794 13568
rect 32866 13496 32898 13568
rect 32498 13484 32898 13496
rect 3698 12480 4098 12492
rect 3698 12408 3730 12480
rect 3802 12408 3818 12480
rect 3890 12408 3906 12480
rect 3978 12408 3994 12480
rect 4066 12408 4098 12480
rect 3698 12396 4098 12408
rect 98 11937 498 11948
rect 98 11864 130 11937
rect 202 11864 218 11937
rect 290 11864 306 11937
rect 378 11864 394 11937
rect 466 11864 498 11937
rect 98 11852 498 11864
rect 3698 11392 4098 11404
rect 3698 11320 3730 11392
rect 3802 11320 3818 11392
rect 3890 11320 3906 11392
rect 3978 11320 3994 11392
rect 4066 11320 4098 11392
rect 3698 11308 4098 11320
rect 10898 11392 11298 11404
rect 10898 11320 10930 11392
rect 11002 11320 11018 11392
rect 11090 11320 11106 11392
rect 11178 11320 11194 11392
rect 11266 11320 11298 11392
rect 10898 11308 11298 11320
rect 18098 11392 18498 11404
rect 18098 11320 18130 11392
rect 18202 11320 18218 11392
rect 18290 11320 18306 11392
rect 18378 11320 18394 11392
rect 18466 11320 18498 11392
rect 18098 11308 18498 11320
rect 25298 11392 25698 11404
rect 25298 11320 25330 11392
rect 25402 11320 25418 11392
rect 25490 11320 25506 11392
rect 25578 11320 25594 11392
rect 25666 11320 25698 11392
rect 25298 11308 25698 11320
rect 32498 11392 32898 11404
rect 32498 11319 32530 11392
rect 32602 11319 32618 11392
rect 32690 11319 32706 11392
rect 32778 11319 32794 11392
rect 32866 11319 32898 11392
rect 32498 11307 32898 11319
rect 3698 9217 4098 9228
rect 3698 9144 3730 9217
rect 3802 9144 3818 9217
rect 3890 9144 3906 9217
rect 3978 9144 3994 9217
rect 4066 9144 4098 9217
rect 3698 9132 4098 9144
rect 10898 9217 11298 9228
rect 10898 9144 10930 9217
rect 11002 9144 11018 9217
rect 11090 9144 11106 9217
rect 11178 9144 11194 9217
rect 11266 9144 11298 9217
rect 10898 9132 11298 9144
rect 18098 9217 18498 9228
rect 18098 9144 18130 9217
rect 18202 9144 18218 9217
rect 18290 9144 18306 9217
rect 18378 9144 18394 9217
rect 18466 9144 18498 9217
rect 18098 9132 18498 9144
rect 25298 9217 25698 9228
rect 25298 9144 25330 9217
rect 25402 9144 25418 9217
rect 25490 9144 25506 9217
rect 25578 9144 25594 9217
rect 25666 9144 25698 9217
rect 25298 9132 25698 9144
rect 32498 9217 32898 9228
rect 32498 9144 32530 9217
rect 32602 9144 32618 9217
rect 32690 9144 32706 9217
rect 32778 9144 32794 9217
rect 32866 9144 32898 9217
rect 32498 9132 32898 9144
rect 3698 7041 4098 7052
rect 3698 6968 3730 7041
rect 3802 6968 3818 7041
rect 3890 6968 3906 7041
rect 3978 6968 3994 7041
rect 4066 6968 4098 7041
rect 3698 6956 4098 6968
rect 10898 7041 11298 7052
rect 10898 6968 10930 7041
rect 11002 6968 11018 7041
rect 11090 6968 11106 7041
rect 11178 6968 11194 7041
rect 11266 6968 11298 7041
rect 10898 6956 11298 6968
rect 25298 7041 25698 7052
rect 25298 6968 25330 7041
rect 25402 6968 25418 7041
rect 25490 6968 25506 7041
rect 25578 6968 25594 7041
rect 25666 6968 25698 7041
rect 25298 6956 25698 6968
rect 32498 7041 32898 7052
rect 32498 6968 32530 7041
rect 32602 6968 32618 7041
rect 32690 6968 32706 7041
rect 32778 6968 32794 7041
rect 32866 6968 32898 7041
rect 32498 6956 32898 6968
rect 7298 6087 7698 6100
rect 7298 6014 7330 6087
rect 7402 6014 7418 6087
rect 7490 6014 7506 6087
rect 7578 6014 7594 6087
rect 7666 6014 7698 6087
rect 7298 6000 7698 6014
rect 14498 6087 14898 6100
rect 14498 6014 14530 6087
rect 14602 6014 14618 6087
rect 14690 6014 14706 6087
rect 14778 6014 14794 6087
rect 14866 6014 14898 6087
rect 14498 6000 14898 6014
rect 21698 6087 22098 6100
rect 21698 6014 21730 6087
rect 21802 6014 21818 6087
rect 21890 6014 21906 6087
rect 21978 6014 21994 6087
rect 22066 6014 22098 6087
rect 21698 6000 22098 6014
rect 28898 6087 29298 6100
rect 28898 6014 28930 6087
rect 29002 6014 29018 6087
rect 29090 6014 29106 6087
rect 29178 6014 29194 6087
rect 29266 6014 29298 6087
rect 28898 6000 29298 6014
use power_ring_2_2  power_ring_2_2_0
timestamp 1623170494
transform 1 0 -26902 0 1 -3400
box 27000 1800 63400 25600
use ring_osc  ring_osc_0
timestamp 1623172293
transform 1 0 0 0 1 6460
box 0 -258 36700 7874
use pwell_co_ring  pwell_co_ring_0
timestamp 1623122433
transform 1 0 0 0 1 0
box 176 6000 36124 14500
<< labels >>
flabel metal2 29854 6202 30014 6402 1 FreeSans 2400 0 0 0 p[0]
port 1 nsew signal output
flabel metal2 23954 6202 24114 6402 1 FreeSans 2400 0 0 0 p[1]
port 2 nsew signal output
flabel metal2 18054 6202 18214 6402 1 FreeSans 2400 0 0 0 p[2]
port 3 nsew signal output
flabel metal2 12154 6202 12314 6402 1 FreeSans 2400 0 0 0 p[3]
port 4 nsew signal output
flabel metal2 6254 6202 6414 6402 1 FreeSans 2400 0 0 0 p[4]
port 5 nsew signal output
flabel metal2 33272 6202 33432 6402 1 FreeSans 2400 0 0 0 p[10]
port 11 nsew signal output
flabel metal2 9364 14134 9524 14334 1 FreeSans 2400 0 0 0 p[6]
port 7 nsew signal output
flabel metal2 15264 14134 15424 14334 1 FreeSans 2400 0 0 0 p[7]
port 8 nsew signal output
flabel metal2 21164 14134 21324 14334 1 FreeSans 2400 0 0 0 p[8]
port 9 nsew signal output
flabel metal2 27064 14134 27224 14334 1 FreeSans 2400 0 0 0 p[9]
port 10 nsew signal output
flabel locali s 781 12099 873 12245 1 FreeSans 2400 0 0 0 enable
port 15 nsew signal input
flabel locali 1327 12275 1496 12335 1 FreeSans 400 0 0 0 hi_logic
flabel metal1 31002 10762 31520 10860 1 FreeSans 2 0 0 0 v_crt
flabel metal1 9336 12652 9634 12780 1 FreeSans 2 0 0 0 pn[6]
flabel metal1 15248 12654 15546 12782 1 FreeSans 2 0 0 0 pn[7]
flabel metal1 21152 12652 21450 12780 1 FreeSans 2 0 0 0 pn[8]
flabel metal1 27044 12652 27342 12780 1 FreeSans 2 0 0 0 pn[9]
flabel metal1 29768 7754 30066 7882 1 FreeSans 2 0 0 0 pn[0]
flabel metal1 23852 7754 24150 7882 1 FreeSans 2 0 0 0 pn[1]
flabel metal1 17956 7754 18254 7882 1 FreeSans 2 0 0 0 pn[2]
flabel metal1 12044 7754 12342 7882 1 FreeSans 2 0 0 0 pn[3]
flabel metal1 6144 7756 6442 7884 1 FreeSans 2 0 0 0 pn[4]
flabel metal2 800 10332 1116 10470 1 FreeSans 2 0 0 0 pn[5]
flabel metal2 34364 9848 34680 9986 1 FreeSans 2 0 0 0 pn[10]
flabel locali 1786 12216 1830 12260 1 FreeSans 2 0 0 0 lo_logic
flabel metal2 2654 6202 2814 6402 1 FreeSans 2400 0 0 0 p[5]
port 6 nsew signal output
flabel locali 954 12118 978 12144 1 FreeSans 300 0 0 0 net3
flabel pdiff 1052 12300 1084 12334 1 FreeSans 300 0 0 0 net1
flabel ndiff 1054 11992 1082 12024 1 FreeSans 300 0 0 0 net2
flabel metal2 36500 10748 36700 10908 1 FreeSans 2400 0 0 0 input_analog
port 12 nsew signal input
flabel metal3 s 30800 21800 31800 22200 1 FreeSans 2400 0 0 0 vccd2
port 13 nsew power bidirectional abutment
flabel metal3 s 30800 20600 31800 21000 1 FreeSans 2400 0 0 0 vssd2
port 14 nsew ground bidirectional abutment
<< end >>
