magic
tech sky130A
timestamp 1637401559
<< psubdiff >>
rect 550 3630 590 3660
rect 620 3630 650 3660
rect 680 3630 710 3660
rect 740 3630 770 3660
rect 800 3630 830 3660
rect 860 3630 890 3660
rect 920 3630 950 3660
rect 980 3630 1010 3660
rect 1040 3630 1070 3660
rect 1100 3630 1130 3660
rect 1160 3630 1190 3660
rect 1220 3630 1250 3660
rect 1280 3630 1310 3660
rect 1340 3630 1370 3660
rect 1400 3630 1430 3660
rect 1460 3630 1490 3660
rect 1520 3630 1550 3660
rect 1580 3630 1610 3660
rect 1640 3630 1670 3660
rect 1700 3630 1730 3660
rect 1760 3630 1790 3660
rect 1820 3630 1850 3660
rect 1880 3630 1910 3660
rect 1940 3630 1970 3660
rect 2000 3630 2030 3660
rect 2060 3630 2090 3660
rect 2120 3630 2150 3660
rect 2180 3630 2210 3660
rect 2240 3630 2270 3660
rect 2300 3630 2330 3660
rect 2360 3630 2390 3660
rect 2420 3630 2450 3660
rect 2480 3630 2510 3660
rect 2540 3630 2570 3660
rect 2600 3630 2630 3660
rect 2660 3630 2690 3660
rect 2720 3630 2750 3660
rect 2780 3630 2810 3660
rect 2840 3630 2870 3660
rect 2900 3630 2930 3660
rect 2960 3630 2990 3660
rect 3020 3630 3050 3660
rect 3080 3630 3110 3660
rect 3140 3630 3170 3660
rect 3200 3630 3230 3660
rect 3260 3630 3290 3660
rect 3320 3630 3350 3660
rect 3380 3630 3410 3660
rect 3440 3630 3470 3660
rect 3500 3630 3530 3660
rect 3560 3630 3590 3660
rect 3620 3630 3650 3660
rect 3680 3630 3710 3660
rect 3740 3630 3770 3660
rect 3800 3630 3830 3660
rect 3860 3630 3890 3660
rect 3920 3630 3950 3660
rect 3980 3630 4010 3660
rect 4040 3630 4070 3660
rect 4100 3630 4130 3660
rect 4160 3630 4190 3660
rect 4220 3630 4250 3660
rect 4280 3630 4310 3660
rect 4340 3630 4370 3660
rect 4400 3630 4430 3660
rect 4460 3630 4490 3660
rect 4520 3630 4550 3660
rect 4580 3630 4610 3660
rect 4640 3630 4670 3660
rect 4700 3630 4730 3660
rect 4760 3630 4790 3660
rect 4820 3630 4850 3660
rect 4880 3630 4910 3660
rect 4940 3630 4970 3660
rect 5000 3630 5030 3660
rect 5060 3630 5090 3660
rect 5120 3630 5150 3660
rect 5180 3630 5210 3660
rect 5240 3630 5270 3660
rect 5300 3630 5330 3660
rect 5360 3630 5390 3660
rect 5420 3630 5450 3660
rect 5480 3630 5510 3660
rect 5540 3630 5570 3660
rect 5600 3630 5630 3660
rect 5660 3630 5690 3660
rect 5720 3630 5750 3660
rect 5780 3630 5810 3660
rect 5840 3630 5870 3660
rect 5900 3630 5930 3660
rect 5960 3630 5990 3660
rect 6020 3630 6050 3660
rect 6080 3630 6110 3660
rect 6140 3630 6170 3660
rect 6200 3630 6230 3660
rect 6260 3630 6290 3660
rect 6320 3630 6350 3660
rect 6380 3630 6410 3660
rect 6440 3630 6470 3660
rect 6500 3630 6530 3660
rect 6560 3630 6590 3660
rect 6620 3630 6650 3660
rect 6680 3630 6710 3660
rect 6740 3630 6770 3660
rect 6800 3630 6830 3660
rect 6860 3630 6890 3660
rect 6920 3630 6950 3660
rect 6980 3630 7010 3660
rect 7040 3630 7070 3660
rect 7100 3630 7130 3660
rect 7160 3630 7190 3660
rect 7220 3630 7250 3660
rect 7280 3630 7310 3660
rect 7340 3630 7370 3660
rect 7400 3630 7430 3660
rect 7460 3630 7490 3660
rect 7520 3630 7550 3660
rect 7580 3630 7610 3660
rect 7640 3630 7670 3660
rect 7700 3630 7730 3660
rect 7760 3630 7790 3660
rect 7820 3630 7850 3660
rect 7880 3630 7910 3660
rect 7940 3630 7970 3660
rect 8000 3630 8030 3660
rect 8060 3630 8090 3660
rect 8120 3630 8150 3660
rect 8180 3630 8210 3660
rect 8240 3630 8270 3660
rect 8300 3630 8330 3660
rect 8360 3630 8390 3660
rect 8420 3630 8450 3660
rect 8480 3630 8510 3660
rect 8540 3630 8570 3660
rect 8600 3630 8630 3660
rect 8660 3630 8690 3660
rect 8720 3630 8750 3660
rect 8780 3630 8810 3660
rect 8840 3630 8870 3660
rect 8900 3630 8930 3660
rect 8960 3630 8990 3660
rect 9020 3630 9050 3660
rect 9080 3630 9110 3660
rect 9140 3630 9170 3660
rect 9200 3630 9230 3660
rect 9260 3630 9290 3660
rect 9320 3630 9350 3660
rect 550 3610 580 3630
rect 550 3550 580 3580
rect 550 3490 580 3520
rect 550 3430 580 3460
rect 550 3370 580 3400
rect 550 3310 580 3340
rect 550 3250 580 3280
rect 550 3190 580 3220
rect 550 3130 580 3160
rect 550 3070 580 3100
rect 550 3010 580 3040
rect 550 2950 580 2980
rect 550 2890 580 2920
rect 550 2830 580 2860
rect 550 2770 580 2800
rect 550 2710 580 2740
rect 550 2650 580 2680
rect 550 2590 580 2620
rect 550 2530 580 2560
rect 550 2470 580 2500
rect 550 2410 580 2440
rect 550 2350 580 2380
rect 550 2290 580 2320
rect 550 2230 580 2260
rect 550 2170 580 2200
rect 550 2120 580 2140
rect 550 2060 580 2080
rect 550 2000 580 2020
rect 550 1940 580 1960
rect 550 1845 580 1910
rect 9380 3610 9410 3660
rect 9380 3550 9410 3580
rect 9380 3490 9410 3520
rect 9380 3430 9410 3460
rect 9380 3370 9410 3400
rect 9380 3310 9410 3340
rect 9380 3250 9410 3280
rect 9380 3190 9410 3220
rect 9380 3130 9410 3160
rect 9380 3070 9410 3100
rect 9380 3010 9410 3040
rect 9380 2950 9410 2980
rect 9380 2890 9410 2920
rect 9380 2830 9410 2860
rect 9380 2770 9410 2800
rect 9380 2710 9410 2740
rect 9380 2650 9410 2680
rect 9380 2590 9410 2620
rect 9380 2530 9410 2560
rect 9380 2470 9410 2500
rect 9380 2410 9410 2440
rect 9380 2350 9410 2380
rect 9380 2290 9410 2320
rect 9380 2230 9410 2260
rect 9380 2170 9410 2200
rect 9380 2120 9410 2140
rect 9380 2060 9410 2080
rect 9380 2000 9410 2020
rect 9380 1940 9410 1960
rect 9380 1845 9410 1910
rect 0 1787 30 1845
rect 60 1815 90 1845
rect 120 1815 150 1845
rect 180 1815 210 1845
rect 240 1815 270 1845
rect 300 1815 330 1845
rect 360 1815 390 1845
rect 420 1815 450 1845
rect 480 1815 510 1845
rect 540 1815 570 1845
rect 600 1815 630 1845
rect 660 1815 690 1845
rect 720 1815 740 1845
rect 770 1815 800 1845
rect 830 1815 860 1845
rect 890 1815 920 1845
rect 950 1815 980 1845
rect 1010 1815 1040 1845
rect 1070 1815 1100 1845
rect 1130 1815 1160 1845
rect 1190 1815 1220 1845
rect 1250 1815 1280 1845
rect 1310 1815 1340 1845
rect 1370 1815 1400 1845
rect 1430 1815 1460 1845
rect 1490 1815 1520 1845
rect 1550 1815 1580 1845
rect 1610 1815 1640 1845
rect 1670 1815 1700 1845
rect 1730 1815 1760 1845
rect 1790 1815 1820 1845
rect 1850 1815 1880 1845
rect 1910 1815 1940 1845
rect 1970 1815 2000 1845
rect 2030 1815 2060 1845
rect 2090 1815 2120 1845
rect 2150 1815 2180 1845
rect 2210 1815 2240 1845
rect 2270 1815 2300 1845
rect 2330 1815 2360 1845
rect 2390 1815 2420 1845
rect 2450 1815 2480 1845
rect 2510 1815 2540 1845
rect 2570 1815 2600 1845
rect 2630 1815 2660 1845
rect 2690 1815 2720 1845
rect 2750 1815 2780 1845
rect 2810 1815 2840 1845
rect 2870 1815 2900 1845
rect 2930 1815 2960 1845
rect 2990 1815 3020 1845
rect 3050 1815 3080 1845
rect 3110 1815 3140 1845
rect 3170 1815 3200 1845
rect 3230 1815 3260 1845
rect 3290 1815 3320 1845
rect 3350 1815 3380 1845
rect 3410 1815 3440 1845
rect 3470 1815 3500 1845
rect 3530 1815 3560 1845
rect 3590 1815 3620 1845
rect 3650 1815 3680 1845
rect 3710 1815 3740 1845
rect 3770 1815 3800 1845
rect 3830 1815 3860 1845
rect 3890 1815 3920 1845
rect 3950 1815 3980 1845
rect 4010 1815 4040 1845
rect 4070 1815 4100 1845
rect 4130 1815 4160 1845
rect 4190 1815 4220 1845
rect 4250 1815 4280 1845
rect 4310 1815 4340 1845
rect 4370 1815 4400 1845
rect 4430 1815 4460 1845
rect 4490 1815 4520 1845
rect 4550 1815 4580 1845
rect 4610 1815 4640 1845
rect 4670 1815 4700 1845
rect 4730 1815 4760 1845
rect 4790 1815 4820 1845
rect 4850 1815 4880 1845
rect 4910 1815 4940 1845
rect 4970 1815 5000 1845
rect 5030 1815 5060 1845
rect 5090 1815 5120 1845
rect 5150 1815 5180 1845
rect 5210 1815 5240 1845
rect 5270 1815 5300 1845
rect 5330 1815 5360 1845
rect 5390 1815 5420 1845
rect 5450 1815 5480 1845
rect 5510 1815 5540 1845
rect 5570 1815 5600 1845
rect 5630 1815 5660 1845
rect 5690 1815 5720 1845
rect 5750 1815 5780 1845
rect 5810 1815 5840 1845
rect 5870 1815 5900 1845
rect 5930 1815 5960 1845
rect 5990 1815 6020 1845
rect 6050 1815 6080 1845
rect 6110 1815 6140 1845
rect 6170 1815 6200 1845
rect 6230 1815 6260 1845
rect 6290 1815 6320 1845
rect 6350 1815 6380 1845
rect 6410 1815 6440 1845
rect 6470 1815 6500 1845
rect 6530 1815 6560 1845
rect 6590 1815 6620 1845
rect 6650 1815 6680 1845
rect 6710 1815 6740 1845
rect 6770 1815 6800 1845
rect 6830 1815 6860 1845
rect 6890 1815 6920 1845
rect 6950 1815 6980 1845
rect 7010 1815 7040 1845
rect 7070 1815 7100 1845
rect 7130 1815 7160 1845
rect 7190 1815 7220 1845
rect 7250 1815 7280 1845
rect 7310 1815 7340 1845
rect 7370 1815 7400 1845
rect 7430 1815 7460 1845
rect 7490 1815 7520 1845
rect 7550 1815 7580 1845
rect 7610 1815 7640 1845
rect 7670 1815 7700 1845
rect 7730 1815 7760 1845
rect 7790 1815 7820 1845
rect 7850 1815 7880 1845
rect 7910 1815 7940 1845
rect 7970 1815 8000 1845
rect 8030 1815 8060 1845
rect 8090 1815 8120 1845
rect 8150 1815 8180 1845
rect 8210 1815 8240 1845
rect 8270 1815 8300 1845
rect 8330 1815 8360 1845
rect 8390 1815 8420 1845
rect 8450 1815 8480 1845
rect 8510 1815 8540 1845
rect 8570 1815 8600 1845
rect 8630 1815 8660 1845
rect 8690 1815 8720 1845
rect 8750 1815 8780 1845
rect 8810 1815 8840 1845
rect 8870 1815 8900 1845
rect 8930 1815 8960 1845
rect 8990 1815 9020 1845
rect 9050 1815 9080 1845
rect 9110 1815 9140 1845
rect 9170 1815 9200 1845
rect 9230 1815 9260 1845
rect 9290 1815 9320 1845
rect 9350 1815 9380 1845
rect 9410 1815 9440 1845
rect 9470 1815 9500 1845
rect 9530 1815 9560 1845
rect 9590 1815 9620 1845
rect 9650 1815 9680 1845
rect 9710 1815 9740 1845
rect 9770 1815 9800 1845
rect 9830 1815 9860 1845
rect 9890 1815 9920 1845
rect 9950 1815 9980 1845
rect 10010 1815 10040 1845
rect 10070 1815 10100 1845
rect 10130 1815 10160 1845
rect 10190 1815 10220 1845
rect 10250 1815 10280 1845
rect 10310 1815 10340 1845
rect 10370 1815 10400 1845
rect 10430 1815 10460 1845
rect 10490 1815 10518 1845
rect 10548 1815 10560 1845
rect 0 1727 30 1757
rect 0 1667 30 1697
rect 0 1607 30 1637
rect 0 1547 30 1577
rect 0 1487 30 1517
rect 0 1427 30 1457
rect 0 1367 30 1397
rect 0 1307 30 1337
rect 0 1247 30 1277
rect 0 1187 30 1217
rect 0 1127 30 1157
rect 0 1067 30 1097
rect 0 1007 30 1037
rect 0 947 30 977
rect 0 887 30 917
rect 0 827 30 857
rect 0 767 30 797
rect 0 707 30 737
rect 0 647 30 677
rect 0 587 30 617
rect 0 527 30 557
rect 0 467 30 497
rect 0 407 30 437
rect 0 347 30 377
rect 0 290 30 317
rect 0 230 30 260
rect 0 170 30 200
rect 0 113 30 140
rect 0 30 30 83
rect 10530 1787 10560 1815
rect 10530 1727 10560 1757
rect 10530 1667 10560 1697
rect 10530 1607 10560 1637
rect 10530 1547 10560 1577
rect 10530 1487 10560 1517
rect 10530 1427 10560 1457
rect 10530 1367 10560 1397
rect 10530 1307 10560 1337
rect 10530 1247 10560 1277
rect 10530 1187 10560 1217
rect 10530 1127 10560 1157
rect 10530 1067 10560 1097
rect 10530 1007 10560 1037
rect 10530 947 10560 977
rect 10530 887 10560 917
rect 10530 827 10560 857
rect 10530 767 10560 797
rect 10530 707 10560 737
rect 10530 647 10560 677
rect 10530 587 10560 617
rect 10530 527 10560 557
rect 10530 467 10560 497
rect 10530 407 10560 437
rect 10530 347 10560 377
rect 10530 290 10560 317
rect 10530 230 10560 260
rect 10530 170 10560 200
rect 10530 113 10560 140
rect 10530 30 10560 83
rect 0 0 40 30
rect 70 0 100 30
rect 130 0 160 30
rect 190 0 220 30
rect 250 0 280 30
rect 310 0 340 30
rect 370 0 400 30
rect 430 0 460 30
rect 490 0 520 30
rect 550 0 580 30
rect 610 0 640 30
rect 670 0 700 30
rect 730 0 760 30
rect 790 0 820 30
rect 850 0 880 30
rect 910 0 940 30
rect 970 0 1000 30
rect 1030 0 1060 30
rect 1090 0 1120 30
rect 1150 0 1180 30
rect 1210 0 1240 30
rect 1270 0 1300 30
rect 1330 0 1360 30
rect 1390 0 1420 30
rect 1450 0 1480 30
rect 1510 0 1540 30
rect 1570 0 1600 30
rect 1630 0 1660 30
rect 1690 0 1720 30
rect 1750 0 1780 30
rect 1810 0 1840 30
rect 1870 0 1900 30
rect 1930 0 1960 30
rect 1990 0 2020 30
rect 2050 0 2080 30
rect 2110 0 2140 30
rect 2170 0 2200 30
rect 2230 0 2260 30
rect 2290 0 2320 30
rect 2350 0 2380 30
rect 2410 0 2440 30
rect 2470 0 2500 30
rect 2530 0 2560 30
rect 2590 0 2620 30
rect 2650 0 2680 30
rect 2710 0 2740 30
rect 2770 0 2800 30
rect 2830 0 2860 30
rect 2890 0 2920 30
rect 2950 0 2980 30
rect 3010 0 3040 30
rect 3070 0 3100 30
rect 3130 0 3160 30
rect 3190 0 3220 30
rect 3250 0 3280 30
rect 3310 0 3340 30
rect 3370 0 3400 30
rect 3430 0 3460 30
rect 3490 0 3520 30
rect 3550 0 3580 30
rect 3610 0 3640 30
rect 3670 0 3700 30
rect 3730 0 3760 30
rect 3790 0 3820 30
rect 3850 0 3880 30
rect 3910 0 3940 30
rect 3970 0 4000 30
rect 4030 0 4060 30
rect 4090 0 4120 30
rect 4150 0 4180 30
rect 4210 0 4240 30
rect 4270 0 4300 30
rect 4330 0 4360 30
rect 4390 0 4420 30
rect 4450 0 4480 30
rect 4510 0 4540 30
rect 4570 0 4600 30
rect 4630 0 4660 30
rect 4690 0 4720 30
rect 4750 0 4780 30
rect 4810 0 4840 30
rect 4870 0 4900 30
rect 4930 0 4960 30
rect 4990 0 5020 30
rect 5050 0 5080 30
rect 5110 0 5140 30
rect 5170 0 5200 30
rect 5230 0 5260 30
rect 5290 0 5320 30
rect 5350 0 5380 30
rect 5410 0 5440 30
rect 5470 0 5500 30
rect 5530 0 5560 30
rect 5590 0 5620 30
rect 5650 0 5680 30
rect 5710 0 5740 30
rect 5770 0 5800 30
rect 5830 0 5860 30
rect 5890 0 5920 30
rect 5950 0 5980 30
rect 6010 0 6040 30
rect 6070 0 6100 30
rect 6130 0 6160 30
rect 6190 0 6220 30
rect 6250 0 6280 30
rect 6310 0 6340 30
rect 6370 0 6400 30
rect 6430 0 6460 30
rect 6490 0 6520 30
rect 6550 0 6580 30
rect 6610 0 6640 30
rect 6670 0 6700 30
rect 6730 0 6760 30
rect 6790 0 6820 30
rect 6850 0 6880 30
rect 6910 0 6940 30
rect 6970 0 7000 30
rect 7030 0 7060 30
rect 7090 0 7120 30
rect 7150 0 7180 30
rect 7210 0 7240 30
rect 7270 0 7300 30
rect 7330 0 7360 30
rect 7390 0 7420 30
rect 7450 0 7480 30
rect 7510 0 7540 30
rect 7570 0 7600 30
rect 7630 0 7660 30
rect 7690 0 7720 30
rect 7750 0 7780 30
rect 7810 0 7840 30
rect 7870 0 7900 30
rect 7930 0 7960 30
rect 7990 0 8020 30
rect 8050 0 8080 30
rect 8110 0 8140 30
rect 8170 0 8200 30
rect 8230 0 8260 30
rect 8290 0 8320 30
rect 8350 0 8380 30
rect 8410 0 8440 30
rect 8470 0 8500 30
rect 8530 0 8560 30
rect 8590 0 8620 30
rect 8650 0 8680 30
rect 8710 0 8740 30
rect 8770 0 8800 30
rect 8830 0 8860 30
rect 8890 0 8920 30
rect 8950 0 8980 30
rect 9010 0 9040 30
rect 9070 0 9100 30
rect 9130 0 9160 30
rect 9190 0 9220 30
rect 9250 0 9280 30
rect 9310 0 9340 30
rect 9370 0 9400 30
rect 9430 0 9460 30
rect 9490 0 9520 30
rect 9550 0 9580 30
rect 9610 0 9640 30
rect 9670 0 9700 30
rect 9730 0 9760 30
rect 9790 0 9820 30
rect 9850 0 9880 30
rect 9910 0 9940 30
rect 9970 0 10000 30
rect 10030 0 10060 30
rect 10090 0 10120 30
rect 10150 0 10180 30
rect 10210 0 10240 30
rect 10270 0 10300 30
rect 10330 0 10360 30
rect 10390 0 10420 30
rect 10450 0 10480 30
rect 10510 0 10560 30
<< psubdiffcont >>
rect 590 3630 620 3660
rect 650 3630 680 3660
rect 710 3630 740 3660
rect 770 3630 800 3660
rect 830 3630 860 3660
rect 890 3630 920 3660
rect 950 3630 980 3660
rect 1010 3630 1040 3660
rect 1070 3630 1100 3660
rect 1130 3630 1160 3660
rect 1190 3630 1220 3660
rect 1250 3630 1280 3660
rect 1310 3630 1340 3660
rect 1370 3630 1400 3660
rect 1430 3630 1460 3660
rect 1490 3630 1520 3660
rect 1550 3630 1580 3660
rect 1610 3630 1640 3660
rect 1670 3630 1700 3660
rect 1730 3630 1760 3660
rect 1790 3630 1820 3660
rect 1850 3630 1880 3660
rect 1910 3630 1940 3660
rect 1970 3630 2000 3660
rect 2030 3630 2060 3660
rect 2090 3630 2120 3660
rect 2150 3630 2180 3660
rect 2210 3630 2240 3660
rect 2270 3630 2300 3660
rect 2330 3630 2360 3660
rect 2390 3630 2420 3660
rect 2450 3630 2480 3660
rect 2510 3630 2540 3660
rect 2570 3630 2600 3660
rect 2630 3630 2660 3660
rect 2690 3630 2720 3660
rect 2750 3630 2780 3660
rect 2810 3630 2840 3660
rect 2870 3630 2900 3660
rect 2930 3630 2960 3660
rect 2990 3630 3020 3660
rect 3050 3630 3080 3660
rect 3110 3630 3140 3660
rect 3170 3630 3200 3660
rect 3230 3630 3260 3660
rect 3290 3630 3320 3660
rect 3350 3630 3380 3660
rect 3410 3630 3440 3660
rect 3470 3630 3500 3660
rect 3530 3630 3560 3660
rect 3590 3630 3620 3660
rect 3650 3630 3680 3660
rect 3710 3630 3740 3660
rect 3770 3630 3800 3660
rect 3830 3630 3860 3660
rect 3890 3630 3920 3660
rect 3950 3630 3980 3660
rect 4010 3630 4040 3660
rect 4070 3630 4100 3660
rect 4130 3630 4160 3660
rect 4190 3630 4220 3660
rect 4250 3630 4280 3660
rect 4310 3630 4340 3660
rect 4370 3630 4400 3660
rect 4430 3630 4460 3660
rect 4490 3630 4520 3660
rect 4550 3630 4580 3660
rect 4610 3630 4640 3660
rect 4670 3630 4700 3660
rect 4730 3630 4760 3660
rect 4790 3630 4820 3660
rect 4850 3630 4880 3660
rect 4910 3630 4940 3660
rect 4970 3630 5000 3660
rect 5030 3630 5060 3660
rect 5090 3630 5120 3660
rect 5150 3630 5180 3660
rect 5210 3630 5240 3660
rect 5270 3630 5300 3660
rect 5330 3630 5360 3660
rect 5390 3630 5420 3660
rect 5450 3630 5480 3660
rect 5510 3630 5540 3660
rect 5570 3630 5600 3660
rect 5630 3630 5660 3660
rect 5690 3630 5720 3660
rect 5750 3630 5780 3660
rect 5810 3630 5840 3660
rect 5870 3630 5900 3660
rect 5930 3630 5960 3660
rect 5990 3630 6020 3660
rect 6050 3630 6080 3660
rect 6110 3630 6140 3660
rect 6170 3630 6200 3660
rect 6230 3630 6260 3660
rect 6290 3630 6320 3660
rect 6350 3630 6380 3660
rect 6410 3630 6440 3660
rect 6470 3630 6500 3660
rect 6530 3630 6560 3660
rect 6590 3630 6620 3660
rect 6650 3630 6680 3660
rect 6710 3630 6740 3660
rect 6770 3630 6800 3660
rect 6830 3630 6860 3660
rect 6890 3630 6920 3660
rect 6950 3630 6980 3660
rect 7010 3630 7040 3660
rect 7070 3630 7100 3660
rect 7130 3630 7160 3660
rect 7190 3630 7220 3660
rect 7250 3630 7280 3660
rect 7310 3630 7340 3660
rect 7370 3630 7400 3660
rect 7430 3630 7460 3660
rect 7490 3630 7520 3660
rect 7550 3630 7580 3660
rect 7610 3630 7640 3660
rect 7670 3630 7700 3660
rect 7730 3630 7760 3660
rect 7790 3630 7820 3660
rect 7850 3630 7880 3660
rect 7910 3630 7940 3660
rect 7970 3630 8000 3660
rect 8030 3630 8060 3660
rect 8090 3630 8120 3660
rect 8150 3630 8180 3660
rect 8210 3630 8240 3660
rect 8270 3630 8300 3660
rect 8330 3630 8360 3660
rect 8390 3630 8420 3660
rect 8450 3630 8480 3660
rect 8510 3630 8540 3660
rect 8570 3630 8600 3660
rect 8630 3630 8660 3660
rect 8690 3630 8720 3660
rect 8750 3630 8780 3660
rect 8810 3630 8840 3660
rect 8870 3630 8900 3660
rect 8930 3630 8960 3660
rect 8990 3630 9020 3660
rect 9050 3630 9080 3660
rect 9110 3630 9140 3660
rect 9170 3630 9200 3660
rect 9230 3630 9260 3660
rect 9290 3630 9320 3660
rect 9350 3630 9380 3660
rect 550 3580 580 3610
rect 550 3520 580 3550
rect 550 3460 580 3490
rect 550 3400 580 3430
rect 550 3340 580 3370
rect 550 3280 580 3310
rect 550 3220 580 3250
rect 550 3160 580 3190
rect 550 3100 580 3130
rect 550 3040 580 3070
rect 550 2980 580 3010
rect 550 2920 580 2950
rect 550 2860 580 2890
rect 550 2800 580 2830
rect 550 2740 580 2770
rect 550 2680 580 2710
rect 550 2620 580 2650
rect 550 2560 580 2590
rect 550 2500 580 2530
rect 550 2440 580 2470
rect 550 2380 580 2410
rect 550 2320 580 2350
rect 550 2260 580 2290
rect 550 2200 580 2230
rect 550 2140 580 2170
rect 550 2080 580 2120
rect 550 2020 580 2060
rect 550 1960 580 2000
rect 550 1910 580 1940
rect 9380 3580 9410 3610
rect 9380 3520 9410 3550
rect 9380 3460 9410 3490
rect 9380 3400 9410 3430
rect 9380 3340 9410 3370
rect 9380 3280 9410 3310
rect 9380 3220 9410 3250
rect 9380 3160 9410 3190
rect 9380 3100 9410 3130
rect 9380 3040 9410 3070
rect 9380 2980 9410 3010
rect 9380 2920 9410 2950
rect 9380 2860 9410 2890
rect 9380 2800 9410 2830
rect 9380 2740 9410 2770
rect 9380 2680 9410 2710
rect 9380 2620 9410 2650
rect 9380 2560 9410 2590
rect 9380 2500 9410 2530
rect 9380 2440 9410 2470
rect 9380 2380 9410 2410
rect 9380 2320 9410 2350
rect 9380 2260 9410 2290
rect 9380 2200 9410 2230
rect 9380 2140 9410 2170
rect 9380 2080 9410 2120
rect 9380 2020 9410 2060
rect 9380 1960 9410 2000
rect 9380 1910 9410 1940
rect 30 1815 60 1845
rect 90 1815 120 1845
rect 150 1815 180 1845
rect 210 1815 240 1845
rect 270 1815 300 1845
rect 330 1815 360 1845
rect 390 1815 420 1845
rect 450 1815 480 1845
rect 510 1815 540 1845
rect 570 1815 600 1845
rect 630 1815 660 1845
rect 690 1815 720 1845
rect 740 1815 770 1845
rect 800 1815 830 1845
rect 860 1815 890 1845
rect 920 1815 950 1845
rect 980 1815 1010 1845
rect 1040 1815 1070 1845
rect 1100 1815 1130 1845
rect 1160 1815 1190 1845
rect 1220 1815 1250 1845
rect 1280 1815 1310 1845
rect 1340 1815 1370 1845
rect 1400 1815 1430 1845
rect 1460 1815 1490 1845
rect 1520 1815 1550 1845
rect 1580 1815 1610 1845
rect 1640 1815 1670 1845
rect 1700 1815 1730 1845
rect 1760 1815 1790 1845
rect 1820 1815 1850 1845
rect 1880 1815 1910 1845
rect 1940 1815 1970 1845
rect 2000 1815 2030 1845
rect 2060 1815 2090 1845
rect 2120 1815 2150 1845
rect 2180 1815 2210 1845
rect 2240 1815 2270 1845
rect 2300 1815 2330 1845
rect 2360 1815 2390 1845
rect 2420 1815 2450 1845
rect 2480 1815 2510 1845
rect 2540 1815 2570 1845
rect 2600 1815 2630 1845
rect 2660 1815 2690 1845
rect 2720 1815 2750 1845
rect 2780 1815 2810 1845
rect 2840 1815 2870 1845
rect 2900 1815 2930 1845
rect 2960 1815 2990 1845
rect 3020 1815 3050 1845
rect 3080 1815 3110 1845
rect 3140 1815 3170 1845
rect 3200 1815 3230 1845
rect 3260 1815 3290 1845
rect 3320 1815 3350 1845
rect 3380 1815 3410 1845
rect 3440 1815 3470 1845
rect 3500 1815 3530 1845
rect 3560 1815 3590 1845
rect 3620 1815 3650 1845
rect 3680 1815 3710 1845
rect 3740 1815 3770 1845
rect 3800 1815 3830 1845
rect 3860 1815 3890 1845
rect 3920 1815 3950 1845
rect 3980 1815 4010 1845
rect 4040 1815 4070 1845
rect 4100 1815 4130 1845
rect 4160 1815 4190 1845
rect 4220 1815 4250 1845
rect 4280 1815 4310 1845
rect 4340 1815 4370 1845
rect 4400 1815 4430 1845
rect 4460 1815 4490 1845
rect 4520 1815 4550 1845
rect 4580 1815 4610 1845
rect 4640 1815 4670 1845
rect 4700 1815 4730 1845
rect 4760 1815 4790 1845
rect 4820 1815 4850 1845
rect 4880 1815 4910 1845
rect 4940 1815 4970 1845
rect 5000 1815 5030 1845
rect 5060 1815 5090 1845
rect 5120 1815 5150 1845
rect 5180 1815 5210 1845
rect 5240 1815 5270 1845
rect 5300 1815 5330 1845
rect 5360 1815 5390 1845
rect 5420 1815 5450 1845
rect 5480 1815 5510 1845
rect 5540 1815 5570 1845
rect 5600 1815 5630 1845
rect 5660 1815 5690 1845
rect 5720 1815 5750 1845
rect 5780 1815 5810 1845
rect 5840 1815 5870 1845
rect 5900 1815 5930 1845
rect 5960 1815 5990 1845
rect 6020 1815 6050 1845
rect 6080 1815 6110 1845
rect 6140 1815 6170 1845
rect 6200 1815 6230 1845
rect 6260 1815 6290 1845
rect 6320 1815 6350 1845
rect 6380 1815 6410 1845
rect 6440 1815 6470 1845
rect 6500 1815 6530 1845
rect 6560 1815 6590 1845
rect 6620 1815 6650 1845
rect 6680 1815 6710 1845
rect 6740 1815 6770 1845
rect 6800 1815 6830 1845
rect 6860 1815 6890 1845
rect 6920 1815 6950 1845
rect 6980 1815 7010 1845
rect 7040 1815 7070 1845
rect 7100 1815 7130 1845
rect 7160 1815 7190 1845
rect 7220 1815 7250 1845
rect 7280 1815 7310 1845
rect 7340 1815 7370 1845
rect 7400 1815 7430 1845
rect 7460 1815 7490 1845
rect 7520 1815 7550 1845
rect 7580 1815 7610 1845
rect 7640 1815 7670 1845
rect 7700 1815 7730 1845
rect 7760 1815 7790 1845
rect 7820 1815 7850 1845
rect 7880 1815 7910 1845
rect 7940 1815 7970 1845
rect 8000 1815 8030 1845
rect 8060 1815 8090 1845
rect 8120 1815 8150 1845
rect 8180 1815 8210 1845
rect 8240 1815 8270 1845
rect 8300 1815 8330 1845
rect 8360 1815 8390 1845
rect 8420 1815 8450 1845
rect 8480 1815 8510 1845
rect 8540 1815 8570 1845
rect 8600 1815 8630 1845
rect 8660 1815 8690 1845
rect 8720 1815 8750 1845
rect 8780 1815 8810 1845
rect 8840 1815 8870 1845
rect 8900 1815 8930 1845
rect 8960 1815 8990 1845
rect 9020 1815 9050 1845
rect 9080 1815 9110 1845
rect 9140 1815 9170 1845
rect 9200 1815 9230 1845
rect 9260 1815 9290 1845
rect 9320 1815 9350 1845
rect 9380 1815 9410 1845
rect 9440 1815 9470 1845
rect 9500 1815 9530 1845
rect 9560 1815 9590 1845
rect 9620 1815 9650 1845
rect 9680 1815 9710 1845
rect 9740 1815 9770 1845
rect 9800 1815 9830 1845
rect 9860 1815 9890 1845
rect 9920 1815 9950 1845
rect 9980 1815 10010 1845
rect 10040 1815 10070 1845
rect 10100 1815 10130 1845
rect 10160 1815 10190 1845
rect 10220 1815 10250 1845
rect 10280 1815 10310 1845
rect 10340 1815 10370 1845
rect 10400 1815 10430 1845
rect 10460 1815 10490 1845
rect 10518 1815 10548 1845
rect 0 1757 30 1787
rect 0 1697 30 1727
rect 0 1637 30 1667
rect 0 1577 30 1607
rect 0 1517 30 1547
rect 0 1457 30 1487
rect 0 1397 30 1427
rect 0 1337 30 1367
rect 0 1277 30 1307
rect 0 1217 30 1247
rect 0 1157 30 1187
rect 0 1097 30 1127
rect 0 1037 30 1067
rect 0 977 30 1007
rect 0 917 30 947
rect 0 857 30 887
rect 0 797 30 827
rect 0 737 30 767
rect 0 677 30 707
rect 0 617 30 647
rect 0 557 30 587
rect 0 497 30 527
rect 0 437 30 467
rect 0 377 30 407
rect 0 317 30 347
rect 0 260 30 290
rect 0 200 30 230
rect 0 140 30 170
rect 0 83 30 113
rect 10530 1757 10560 1787
rect 10530 1697 10560 1727
rect 10530 1637 10560 1667
rect 10530 1577 10560 1607
rect 10530 1517 10560 1547
rect 10530 1457 10560 1487
rect 10530 1397 10560 1427
rect 10530 1337 10560 1367
rect 10530 1277 10560 1307
rect 10530 1217 10560 1247
rect 10530 1157 10560 1187
rect 10530 1097 10560 1127
rect 10530 1037 10560 1067
rect 10530 977 10560 1007
rect 10530 917 10560 947
rect 10530 857 10560 887
rect 10530 797 10560 827
rect 10530 737 10560 767
rect 10530 677 10560 707
rect 10530 617 10560 647
rect 10530 557 10560 587
rect 10530 497 10560 527
rect 10530 437 10560 467
rect 10530 377 10560 407
rect 10530 317 10560 347
rect 10530 260 10560 290
rect 10530 200 10560 230
rect 10530 140 10560 170
rect 10530 83 10560 113
rect 40 0 70 30
rect 100 0 130 30
rect 160 0 190 30
rect 220 0 250 30
rect 280 0 310 30
rect 340 0 370 30
rect 400 0 430 30
rect 460 0 490 30
rect 520 0 550 30
rect 580 0 610 30
rect 640 0 670 30
rect 700 0 730 30
rect 760 0 790 30
rect 820 0 850 30
rect 880 0 910 30
rect 940 0 970 30
rect 1000 0 1030 30
rect 1060 0 1090 30
rect 1120 0 1150 30
rect 1180 0 1210 30
rect 1240 0 1270 30
rect 1300 0 1330 30
rect 1360 0 1390 30
rect 1420 0 1450 30
rect 1480 0 1510 30
rect 1540 0 1570 30
rect 1600 0 1630 30
rect 1660 0 1690 30
rect 1720 0 1750 30
rect 1780 0 1810 30
rect 1840 0 1870 30
rect 1900 0 1930 30
rect 1960 0 1990 30
rect 2020 0 2050 30
rect 2080 0 2110 30
rect 2140 0 2170 30
rect 2200 0 2230 30
rect 2260 0 2290 30
rect 2320 0 2350 30
rect 2380 0 2410 30
rect 2440 0 2470 30
rect 2500 0 2530 30
rect 2560 0 2590 30
rect 2620 0 2650 30
rect 2680 0 2710 30
rect 2740 0 2770 30
rect 2800 0 2830 30
rect 2860 0 2890 30
rect 2920 0 2950 30
rect 2980 0 3010 30
rect 3040 0 3070 30
rect 3100 0 3130 30
rect 3160 0 3190 30
rect 3220 0 3250 30
rect 3280 0 3310 30
rect 3340 0 3370 30
rect 3400 0 3430 30
rect 3460 0 3490 30
rect 3520 0 3550 30
rect 3580 0 3610 30
rect 3640 0 3670 30
rect 3700 0 3730 30
rect 3760 0 3790 30
rect 3820 0 3850 30
rect 3880 0 3910 30
rect 3940 0 3970 30
rect 4000 0 4030 30
rect 4060 0 4090 30
rect 4120 0 4150 30
rect 4180 0 4210 30
rect 4240 0 4270 30
rect 4300 0 4330 30
rect 4360 0 4390 30
rect 4420 0 4450 30
rect 4480 0 4510 30
rect 4540 0 4570 30
rect 4600 0 4630 30
rect 4660 0 4690 30
rect 4720 0 4750 30
rect 4780 0 4810 30
rect 4840 0 4870 30
rect 4900 0 4930 30
rect 4960 0 4990 30
rect 5020 0 5050 30
rect 5080 0 5110 30
rect 5140 0 5170 30
rect 5200 0 5230 30
rect 5260 0 5290 30
rect 5320 0 5350 30
rect 5380 0 5410 30
rect 5440 0 5470 30
rect 5500 0 5530 30
rect 5560 0 5590 30
rect 5620 0 5650 30
rect 5680 0 5710 30
rect 5740 0 5770 30
rect 5800 0 5830 30
rect 5860 0 5890 30
rect 5920 0 5950 30
rect 5980 0 6010 30
rect 6040 0 6070 30
rect 6100 0 6130 30
rect 6160 0 6190 30
rect 6220 0 6250 30
rect 6280 0 6310 30
rect 6340 0 6370 30
rect 6400 0 6430 30
rect 6460 0 6490 30
rect 6520 0 6550 30
rect 6580 0 6610 30
rect 6640 0 6670 30
rect 6700 0 6730 30
rect 6760 0 6790 30
rect 6820 0 6850 30
rect 6880 0 6910 30
rect 6940 0 6970 30
rect 7000 0 7030 30
rect 7060 0 7090 30
rect 7120 0 7150 30
rect 7180 0 7210 30
rect 7240 0 7270 30
rect 7300 0 7330 30
rect 7360 0 7390 30
rect 7420 0 7450 30
rect 7480 0 7510 30
rect 7540 0 7570 30
rect 7600 0 7630 30
rect 7660 0 7690 30
rect 7720 0 7750 30
rect 7780 0 7810 30
rect 7840 0 7870 30
rect 7900 0 7930 30
rect 7960 0 7990 30
rect 8020 0 8050 30
rect 8080 0 8110 30
rect 8140 0 8170 30
rect 8200 0 8230 30
rect 8260 0 8290 30
rect 8320 0 8350 30
rect 8380 0 8410 30
rect 8440 0 8470 30
rect 8500 0 8530 30
rect 8560 0 8590 30
rect 8620 0 8650 30
rect 8680 0 8710 30
rect 8740 0 8770 30
rect 8800 0 8830 30
rect 8860 0 8890 30
rect 8920 0 8950 30
rect 8980 0 9010 30
rect 9040 0 9070 30
rect 9100 0 9130 30
rect 9160 0 9190 30
rect 9220 0 9250 30
rect 9280 0 9310 30
rect 9340 0 9370 30
rect 9400 0 9430 30
rect 9460 0 9490 30
rect 9520 0 9550 30
rect 9580 0 9610 30
rect 9640 0 9670 30
rect 9700 0 9730 30
rect 9760 0 9790 30
rect 9820 0 9850 30
rect 9880 0 9910 30
rect 9940 0 9970 30
rect 10000 0 10030 30
rect 10060 0 10090 30
rect 10120 0 10150 30
rect 10180 0 10210 30
rect 10240 0 10270 30
rect 10300 0 10330 30
rect 10360 0 10390 30
rect 10420 0 10450 30
rect 10480 0 10510 30
<< locali >>
rect 550 3630 590 3660
rect 620 3630 650 3660
rect 680 3630 710 3660
rect 740 3630 770 3660
rect 800 3630 830 3660
rect 860 3630 890 3660
rect 920 3630 950 3660
rect 980 3630 1010 3660
rect 1040 3630 1070 3660
rect 1100 3630 1130 3660
rect 1160 3630 1190 3660
rect 1220 3630 1250 3660
rect 1280 3630 1310 3660
rect 1340 3630 1370 3660
rect 1400 3630 1430 3660
rect 1460 3630 1490 3660
rect 1520 3630 1550 3660
rect 1580 3630 1610 3660
rect 1640 3630 1670 3660
rect 1700 3630 1730 3660
rect 1760 3630 1790 3660
rect 1820 3630 1850 3660
rect 1880 3630 1910 3660
rect 1940 3630 1970 3660
rect 2000 3630 2030 3660
rect 2060 3630 2090 3660
rect 2120 3630 2150 3660
rect 2180 3630 2210 3660
rect 2240 3630 2270 3660
rect 2300 3630 2330 3660
rect 2360 3630 2390 3660
rect 2420 3630 2450 3660
rect 2480 3630 2510 3660
rect 2540 3630 2570 3660
rect 2600 3630 2630 3660
rect 2660 3630 2690 3660
rect 2720 3630 2750 3660
rect 2780 3630 2810 3660
rect 2840 3630 2870 3660
rect 2900 3630 2930 3660
rect 2960 3630 2990 3660
rect 3020 3630 3050 3660
rect 3080 3630 3110 3660
rect 3140 3630 3170 3660
rect 3200 3630 3230 3660
rect 3260 3630 3290 3660
rect 3320 3630 3350 3660
rect 3380 3630 3410 3660
rect 3440 3630 3470 3660
rect 3500 3630 3530 3660
rect 3560 3630 3590 3660
rect 3620 3630 3650 3660
rect 3680 3630 3710 3660
rect 3740 3630 3770 3660
rect 3800 3630 3830 3660
rect 3860 3630 3890 3660
rect 3920 3630 3950 3660
rect 3980 3630 4010 3660
rect 4040 3630 4070 3660
rect 4100 3630 4130 3660
rect 4160 3630 4190 3660
rect 4220 3630 4250 3660
rect 4280 3630 4310 3660
rect 4340 3630 4370 3660
rect 4400 3630 4430 3660
rect 4460 3630 4490 3660
rect 4520 3630 4550 3660
rect 4580 3630 4610 3660
rect 4640 3630 4670 3660
rect 4700 3630 4730 3660
rect 4760 3630 4790 3660
rect 4820 3630 4850 3660
rect 4880 3630 4910 3660
rect 4940 3630 4970 3660
rect 5000 3630 5030 3660
rect 5060 3630 5090 3660
rect 5120 3630 5150 3660
rect 5180 3630 5210 3660
rect 5240 3630 5270 3660
rect 5300 3630 5330 3660
rect 5360 3630 5390 3660
rect 5420 3630 5450 3660
rect 5480 3630 5510 3660
rect 5540 3630 5570 3660
rect 5600 3630 5630 3660
rect 5660 3630 5690 3660
rect 5720 3630 5750 3660
rect 5780 3630 5810 3660
rect 5840 3630 5870 3660
rect 5900 3630 5930 3660
rect 5960 3630 5990 3660
rect 6020 3630 6050 3660
rect 6080 3630 6110 3660
rect 6140 3630 6170 3660
rect 6200 3630 6230 3660
rect 6260 3630 6290 3660
rect 6320 3630 6350 3660
rect 6380 3630 6410 3660
rect 6440 3630 6470 3660
rect 6500 3630 6530 3660
rect 6560 3630 6590 3660
rect 6620 3630 6650 3660
rect 6680 3630 6710 3660
rect 6740 3630 6770 3660
rect 6800 3630 6830 3660
rect 6860 3630 6890 3660
rect 6920 3630 6950 3660
rect 6980 3630 7010 3660
rect 7040 3630 7070 3660
rect 7100 3630 7130 3660
rect 7160 3630 7190 3660
rect 7220 3630 7250 3660
rect 7280 3630 7310 3660
rect 7340 3630 7370 3660
rect 7400 3630 7430 3660
rect 7460 3630 7490 3660
rect 7520 3630 7550 3660
rect 7580 3630 7610 3660
rect 7640 3630 7670 3660
rect 7700 3630 7730 3660
rect 7760 3630 7790 3660
rect 7820 3630 7850 3660
rect 7880 3630 7910 3660
rect 7940 3630 7970 3660
rect 8000 3630 8030 3660
rect 8060 3630 8090 3660
rect 8120 3630 8150 3660
rect 8180 3630 8210 3660
rect 8240 3630 8270 3660
rect 8300 3630 8330 3660
rect 8360 3630 8390 3660
rect 8420 3630 8450 3660
rect 8480 3630 8510 3660
rect 8540 3630 8570 3660
rect 8600 3630 8630 3660
rect 8660 3630 8690 3660
rect 8720 3630 8750 3660
rect 8780 3630 8810 3660
rect 8840 3630 8870 3660
rect 8900 3630 8930 3660
rect 8960 3630 8990 3660
rect 9020 3630 9050 3660
rect 9080 3630 9110 3660
rect 9140 3630 9170 3660
rect 9200 3630 9230 3660
rect 9260 3630 9290 3660
rect 9320 3630 9350 3660
rect 550 3610 580 3630
rect 550 3550 580 3580
rect 550 3490 580 3520
rect 550 3430 580 3460
rect 550 3370 580 3400
rect 550 3310 580 3340
rect 550 3250 580 3280
rect 550 3190 580 3220
rect 550 3130 580 3160
rect 550 3070 580 3100
rect 550 3010 580 3040
rect 550 2950 580 2980
rect 550 2890 580 2920
rect 550 2830 580 2860
rect 550 2770 580 2800
rect 550 2710 580 2740
rect 550 2650 580 2680
rect 550 2590 580 2620
rect 550 2530 580 2560
rect 550 2470 580 2500
rect 550 2410 580 2440
rect 550 2350 580 2380
rect 550 2290 580 2320
rect 550 2230 580 2260
rect 550 2170 580 2200
rect 550 2120 580 2140
rect 550 2060 580 2080
rect 550 2000 580 2020
rect 550 1940 580 1960
rect 550 1845 580 1910
rect 9380 3610 9410 3660
rect 9380 3550 9410 3580
rect 9380 3490 9410 3520
rect 9380 3430 9410 3460
rect 9380 3370 9410 3400
rect 9380 3310 9410 3340
rect 9380 3250 9410 3280
rect 9380 3190 9410 3220
rect 9380 3130 9410 3160
rect 9380 3070 9410 3100
rect 9380 3010 9410 3040
rect 9380 2950 9410 2980
rect 9380 2890 9410 2920
rect 9380 2830 9410 2860
rect 9380 2770 9410 2800
rect 9380 2710 9410 2740
rect 9380 2650 9410 2680
rect 9380 2590 9410 2620
rect 9380 2530 9410 2560
rect 9380 2470 9410 2500
rect 9380 2410 9410 2440
rect 9380 2350 9410 2380
rect 9380 2290 9410 2320
rect 9380 2230 9410 2260
rect 9380 2170 9410 2200
rect 9380 2120 9410 2140
rect 9380 2060 9410 2080
rect 9380 2000 9410 2020
rect 9380 1940 9410 1960
rect 9380 1845 9410 1910
rect 0 1787 30 1845
rect 60 1815 90 1845
rect 120 1815 150 1845
rect 180 1815 210 1845
rect 240 1815 270 1845
rect 300 1815 330 1845
rect 360 1815 390 1845
rect 420 1815 450 1845
rect 480 1815 510 1845
rect 540 1815 570 1845
rect 600 1815 630 1845
rect 660 1815 690 1845
rect 720 1815 740 1845
rect 770 1815 800 1845
rect 830 1815 860 1845
rect 890 1815 920 1845
rect 950 1815 980 1845
rect 1010 1815 1040 1845
rect 1070 1815 1100 1845
rect 1130 1815 1160 1845
rect 1190 1815 1220 1845
rect 1250 1815 1280 1845
rect 1310 1815 1340 1845
rect 1370 1815 1400 1845
rect 1430 1815 1460 1845
rect 1490 1815 1520 1845
rect 1550 1815 1580 1845
rect 1610 1815 1640 1845
rect 1670 1815 1700 1845
rect 1730 1815 1760 1845
rect 1790 1815 1820 1845
rect 1850 1815 1880 1845
rect 1910 1815 1940 1845
rect 1970 1815 2000 1845
rect 2030 1815 2060 1845
rect 2090 1815 2120 1845
rect 2150 1815 2180 1845
rect 2210 1815 2240 1845
rect 2270 1815 2300 1845
rect 2330 1815 2360 1845
rect 2390 1815 2420 1845
rect 2450 1815 2480 1845
rect 2510 1815 2540 1845
rect 2570 1815 2600 1845
rect 2630 1815 2660 1845
rect 2690 1815 2720 1845
rect 2750 1815 2780 1845
rect 2810 1815 2840 1845
rect 2870 1815 2900 1845
rect 2930 1815 2960 1845
rect 2990 1815 3020 1845
rect 3050 1815 3080 1845
rect 3110 1815 3140 1845
rect 3170 1815 3200 1845
rect 3230 1815 3260 1845
rect 3290 1815 3320 1845
rect 3350 1815 3380 1845
rect 3410 1815 3440 1845
rect 3470 1815 3500 1845
rect 3530 1815 3560 1845
rect 3590 1815 3620 1845
rect 3650 1815 3680 1845
rect 3710 1815 3740 1845
rect 3770 1815 3800 1845
rect 3830 1815 3860 1845
rect 3890 1815 3920 1845
rect 3950 1815 3980 1845
rect 4010 1815 4040 1845
rect 4070 1815 4100 1845
rect 4130 1815 4160 1845
rect 4190 1815 4220 1845
rect 4250 1815 4280 1845
rect 4310 1815 4340 1845
rect 4370 1815 4400 1845
rect 4430 1815 4460 1845
rect 4490 1815 4520 1845
rect 4550 1815 4580 1845
rect 4610 1815 4640 1845
rect 4670 1815 4700 1845
rect 4730 1815 4760 1845
rect 4790 1815 4820 1845
rect 4850 1815 4880 1845
rect 4910 1815 4940 1845
rect 4970 1815 5000 1845
rect 5030 1815 5060 1845
rect 5090 1815 5120 1845
rect 5150 1815 5180 1845
rect 5210 1815 5240 1845
rect 5270 1815 5300 1845
rect 5330 1815 5360 1845
rect 5390 1815 5420 1845
rect 5450 1815 5480 1845
rect 5510 1815 5540 1845
rect 5570 1815 5600 1845
rect 5630 1815 5660 1845
rect 5690 1815 5720 1845
rect 5750 1815 5780 1845
rect 5810 1815 5840 1845
rect 5870 1815 5900 1845
rect 5930 1815 5960 1845
rect 5990 1815 6020 1845
rect 6050 1815 6080 1845
rect 6110 1815 6140 1845
rect 6170 1815 6200 1845
rect 6230 1815 6260 1845
rect 6290 1815 6320 1845
rect 6350 1815 6380 1845
rect 6410 1815 6440 1845
rect 6470 1815 6500 1845
rect 6530 1815 6560 1845
rect 6590 1815 6620 1845
rect 6650 1815 6680 1845
rect 6710 1815 6740 1845
rect 6770 1815 6800 1845
rect 6830 1815 6860 1845
rect 6890 1815 6920 1845
rect 6950 1815 6980 1845
rect 7010 1815 7040 1845
rect 7070 1815 7100 1845
rect 7130 1815 7160 1845
rect 7190 1815 7220 1845
rect 7250 1815 7280 1845
rect 7310 1815 7340 1845
rect 7370 1815 7400 1845
rect 7430 1815 7460 1845
rect 7490 1815 7520 1845
rect 7550 1815 7580 1845
rect 7610 1815 7640 1845
rect 7670 1815 7700 1845
rect 7730 1815 7760 1845
rect 7790 1815 7820 1845
rect 7850 1815 7880 1845
rect 7910 1815 7940 1845
rect 7970 1815 8000 1845
rect 8030 1815 8060 1845
rect 8090 1815 8120 1845
rect 8150 1815 8180 1845
rect 8210 1815 8240 1845
rect 8270 1815 8300 1845
rect 8330 1815 8360 1845
rect 8390 1815 8420 1845
rect 8450 1815 8480 1845
rect 8510 1815 8540 1845
rect 8570 1815 8600 1845
rect 8630 1815 8660 1845
rect 8690 1815 8720 1845
rect 8750 1815 8780 1845
rect 8810 1815 8840 1845
rect 8870 1815 8900 1845
rect 8930 1815 8960 1845
rect 8990 1815 9020 1845
rect 9050 1815 9080 1845
rect 9110 1815 9140 1845
rect 9170 1815 9200 1845
rect 9230 1815 9260 1845
rect 9290 1815 9320 1845
rect 9350 1815 9380 1845
rect 9410 1815 9440 1845
rect 9470 1815 9500 1845
rect 9530 1815 9560 1845
rect 9590 1815 9620 1845
rect 9650 1815 9680 1845
rect 9710 1815 9740 1845
rect 9770 1815 9800 1845
rect 9830 1815 9860 1845
rect 9890 1815 9920 1845
rect 9950 1815 9980 1845
rect 10010 1815 10040 1845
rect 10070 1815 10100 1845
rect 10130 1815 10160 1845
rect 10190 1815 10220 1845
rect 10250 1815 10280 1845
rect 10310 1815 10340 1845
rect 10370 1815 10400 1845
rect 10430 1815 10460 1845
rect 10490 1815 10518 1845
rect 10548 1815 10560 1845
rect 0 1727 30 1757
rect 0 1667 30 1697
rect 0 1607 30 1637
rect 0 1547 30 1577
rect 0 1487 30 1517
rect 0 1427 30 1457
rect 0 1367 30 1397
rect 0 1307 30 1337
rect 0 1247 30 1277
rect 0 1187 30 1217
rect 0 1127 30 1157
rect 0 1067 30 1097
rect 0 1007 30 1037
rect 0 947 30 977
rect 0 887 30 917
rect 0 827 30 857
rect 0 767 30 797
rect 0 707 30 737
rect 0 647 30 677
rect 0 587 30 617
rect 0 527 30 557
rect 0 467 30 497
rect 0 407 30 437
rect 0 347 30 377
rect 0 290 30 317
rect 0 230 30 260
rect 0 170 30 200
rect 0 113 30 140
rect 0 30 30 83
rect 10530 1787 10560 1815
rect 10530 1727 10560 1757
rect 10530 1667 10560 1697
rect 10530 1607 10560 1637
rect 10530 1547 10560 1577
rect 10530 1487 10560 1517
rect 10530 1427 10560 1457
rect 10530 1367 10560 1397
rect 10530 1307 10560 1337
rect 10530 1247 10560 1277
rect 10530 1187 10560 1217
rect 10530 1127 10560 1157
rect 10530 1067 10560 1097
rect 10530 1007 10560 1037
rect 10530 947 10560 977
rect 10530 887 10560 917
rect 10530 827 10560 857
rect 10530 767 10560 797
rect 10530 707 10560 737
rect 10530 647 10560 677
rect 10530 587 10560 617
rect 10530 527 10560 557
rect 10530 467 10560 497
rect 10530 407 10560 437
rect 10530 347 10560 377
rect 10530 290 10560 317
rect 10530 230 10560 260
rect 10530 170 10560 200
rect 10530 113 10560 140
rect 10530 30 10560 83
rect 0 0 40 30
rect 70 0 100 30
rect 130 0 160 30
rect 190 0 220 30
rect 250 0 280 30
rect 310 0 340 30
rect 370 0 400 30
rect 430 0 460 30
rect 490 0 520 30
rect 550 0 580 30
rect 610 0 640 30
rect 670 0 700 30
rect 730 0 760 30
rect 790 0 820 30
rect 850 0 880 30
rect 910 0 940 30
rect 970 0 1000 30
rect 1030 0 1060 30
rect 1090 0 1120 30
rect 1150 0 1180 30
rect 1210 0 1240 30
rect 1270 0 1300 30
rect 1330 0 1360 30
rect 1390 0 1420 30
rect 1450 0 1480 30
rect 1510 0 1540 30
rect 1570 0 1600 30
rect 1630 0 1660 30
rect 1690 0 1720 30
rect 1750 0 1780 30
rect 1810 0 1840 30
rect 1870 0 1900 30
rect 1930 0 1960 30
rect 1990 0 2020 30
rect 2050 0 2080 30
rect 2110 0 2140 30
rect 2170 0 2200 30
rect 2230 0 2260 30
rect 2290 0 2320 30
rect 2350 0 2380 30
rect 2410 0 2440 30
rect 2470 0 2500 30
rect 2530 0 2560 30
rect 2590 0 2620 30
rect 2650 0 2680 30
rect 2710 0 2740 30
rect 2770 0 2800 30
rect 2830 0 2860 30
rect 2890 0 2920 30
rect 2950 0 2980 30
rect 3010 0 3040 30
rect 3070 0 3100 30
rect 3130 0 3160 30
rect 3190 0 3220 30
rect 3250 0 3280 30
rect 3310 0 3340 30
rect 3370 0 3400 30
rect 3430 0 3460 30
rect 3490 0 3520 30
rect 3550 0 3580 30
rect 3610 0 3640 30
rect 3670 0 3700 30
rect 3730 0 3760 30
rect 3790 0 3820 30
rect 3850 0 3880 30
rect 3910 0 3940 30
rect 3970 0 4000 30
rect 4030 0 4060 30
rect 4090 0 4120 30
rect 4150 0 4180 30
rect 4210 0 4240 30
rect 4270 0 4300 30
rect 4330 0 4360 30
rect 4390 0 4420 30
rect 4450 0 4480 30
rect 4510 0 4540 30
rect 4570 0 4600 30
rect 4630 0 4660 30
rect 4690 0 4720 30
rect 4750 0 4780 30
rect 4810 0 4840 30
rect 4870 0 4900 30
rect 4930 0 4960 30
rect 4990 0 5020 30
rect 5050 0 5080 30
rect 5110 0 5140 30
rect 5170 0 5200 30
rect 5230 0 5260 30
rect 5290 0 5320 30
rect 5350 0 5380 30
rect 5410 0 5440 30
rect 5470 0 5500 30
rect 5530 0 5560 30
rect 5590 0 5620 30
rect 5650 0 5680 30
rect 5710 0 5740 30
rect 5770 0 5800 30
rect 5830 0 5860 30
rect 5890 0 5920 30
rect 5950 0 5980 30
rect 6010 0 6040 30
rect 6070 0 6100 30
rect 6130 0 6160 30
rect 6190 0 6220 30
rect 6250 0 6280 30
rect 6310 0 6340 30
rect 6370 0 6400 30
rect 6430 0 6460 30
rect 6490 0 6520 30
rect 6550 0 6580 30
rect 6610 0 6640 30
rect 6670 0 6700 30
rect 6730 0 6760 30
rect 6790 0 6820 30
rect 6850 0 6880 30
rect 6910 0 6940 30
rect 6970 0 7000 30
rect 7030 0 7060 30
rect 7090 0 7120 30
rect 7150 0 7180 30
rect 7210 0 7240 30
rect 7270 0 7300 30
rect 7330 0 7360 30
rect 7390 0 7420 30
rect 7450 0 7480 30
rect 7510 0 7540 30
rect 7570 0 7600 30
rect 7630 0 7660 30
rect 7690 0 7720 30
rect 7750 0 7780 30
rect 7810 0 7840 30
rect 7870 0 7900 30
rect 7930 0 7960 30
rect 7990 0 8020 30
rect 8050 0 8080 30
rect 8110 0 8140 30
rect 8170 0 8200 30
rect 8230 0 8260 30
rect 8290 0 8320 30
rect 8350 0 8380 30
rect 8410 0 8440 30
rect 8470 0 8500 30
rect 8530 0 8560 30
rect 8590 0 8620 30
rect 8650 0 8680 30
rect 8710 0 8740 30
rect 8770 0 8800 30
rect 8830 0 8860 30
rect 8890 0 8920 30
rect 8950 0 8980 30
rect 9010 0 9040 30
rect 9070 0 9100 30
rect 9130 0 9160 30
rect 9190 0 9220 30
rect 9250 0 9280 30
rect 9310 0 9340 30
rect 9370 0 9400 30
rect 9430 0 9460 30
rect 9490 0 9520 30
rect 9550 0 9580 30
rect 9610 0 9640 30
rect 9670 0 9700 30
rect 9730 0 9760 30
rect 9790 0 9820 30
rect 9850 0 9880 30
rect 9910 0 9940 30
rect 9970 0 10000 30
rect 10030 0 10060 30
rect 10090 0 10120 30
rect 10150 0 10180 30
rect 10210 0 10240 30
rect 10270 0 10300 30
rect 10330 0 10360 30
rect 10390 0 10420 30
rect 10450 0 10480 30
rect 10510 0 10560 30
<< end >>
