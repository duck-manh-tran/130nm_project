magic
tech sky130A
magscale 1 2
timestamp 1623637110
<< pwell >>
rect -400 3308 -328 3380
rect 372 2012 1142 2084
rect 1474 2012 2244 2084
<< poly >>
rect -204 3534 176 3600
rect 234 3534 614 3600
rect -204 3450 614 3534
rect -204 3390 -194 3450
rect -134 3390 -100 3450
rect -40 3390 -6 3450
rect 54 3390 356 3450
rect 416 3390 450 3450
rect 510 3390 544 3450
rect 604 3390 614 3450
rect -204 3314 614 3390
rect -204 3246 176 3314
rect 234 3246 614 3314
rect 900 3534 1280 3600
rect 1338 3534 1718 3600
rect 900 3450 1718 3534
rect 900 3390 910 3450
rect 970 3390 1004 3450
rect 1064 3390 1098 3450
rect 1158 3390 1460 3450
rect 1520 3390 1554 3450
rect 1614 3390 1648 3450
rect 1708 3390 1718 3450
rect 900 3314 1718 3390
rect 900 3246 1280 3314
rect 1338 3246 1718 3314
rect 2004 3450 2384 3582
rect 2004 3390 2014 3450
rect 2074 3390 2108 3450
rect 2168 3390 2202 3450
rect 2262 3390 2384 3450
rect 2004 3258 2384 3390
rect 2670 3450 3050 3582
rect 2670 3390 2680 3450
rect 2740 3390 2774 3450
rect 2834 3390 2868 3450
rect 2928 3390 3050 3450
rect 2670 3258 3050 3390
<< polycont >>
rect -194 3390 -134 3450
rect -100 3390 -40 3450
rect -6 3390 54 3450
rect 356 3390 416 3450
rect 450 3390 510 3450
rect 544 3390 604 3450
rect 910 3390 970 3450
rect 1004 3390 1064 3450
rect 1098 3390 1158 3450
rect 1460 3390 1520 3450
rect 1554 3390 1614 3450
rect 1648 3390 1708 3450
rect 2014 3390 2074 3450
rect 2108 3390 2168 3450
rect 2202 3390 2262 3450
rect 2680 3390 2740 3450
rect 2774 3390 2834 3450
rect 2868 3390 2928 3450
<< locali >>
rect -364 4798 14 4804
rect -364 4738 -352 4798
rect -292 4738 -254 4798
rect -194 4738 -156 4798
rect -96 4738 -58 4798
rect 2 4738 14 4798
rect -364 4732 14 4738
rect 372 4798 1142 4804
rect 372 4738 384 4798
rect 444 4738 482 4798
rect 542 4738 580 4798
rect 640 4738 678 4798
rect 738 4738 776 4798
rect 836 4738 874 4798
rect 934 4738 972 4798
rect 1032 4738 1070 4798
rect 1130 4738 1142 4798
rect 372 4732 1142 4738
rect 1474 4798 2244 4804
rect 1474 4738 1486 4798
rect 1546 4738 1584 4798
rect 1644 4738 1682 4798
rect 1742 4738 1780 4798
rect 1840 4738 1878 4798
rect 1938 4738 1976 4798
rect 2036 4738 2074 4798
rect 2134 4738 2172 4798
rect 2232 4738 2244 4798
rect 1474 4732 2244 4738
rect 2612 4798 2892 4804
rect 2612 4738 2624 4798
rect 2684 4738 2722 4798
rect 2782 4738 2820 4798
rect 2880 4738 2892 4798
rect 2612 4732 2892 4738
rect 175 3722 235 4684
rect -20 3456 56 3466
rect -210 3450 56 3456
rect -134 3390 -112 3450
rect -40 3390 -14 3450
rect 54 3390 56 3450
rect -210 3384 56 3390
rect -20 3374 56 3384
rect -262 2084 -204 3174
rect 175 2166 235 3662
rect 354 3456 430 3466
rect 1084 3456 1160 3466
rect 354 3450 620 3456
rect 354 3390 356 3450
rect 424 3390 450 3450
rect 522 3390 544 3450
rect 354 3384 620 3390
rect 894 3450 1160 3456
rect 970 3390 992 3450
rect 1064 3390 1090 3450
rect 1158 3390 1160 3450
rect 894 3384 1160 3390
rect 354 3374 430 3384
rect 1084 3374 1160 3384
rect 1279 3178 1339 4684
rect 1458 3456 1534 3466
rect 2188 3456 2264 3466
rect 1458 3450 1724 3456
rect 1458 3390 1460 3450
rect 1528 3390 1554 3450
rect 1626 3390 1648 3450
rect 1458 3384 1724 3390
rect 1998 3450 2264 3456
rect 2074 3390 2096 3450
rect 2168 3390 2194 3450
rect 2262 3390 2264 3450
rect 1998 3384 2264 3390
rect 1458 3374 1534 3384
rect 2188 3374 2264 3384
rect 614 2084 672 3174
rect 842 2084 900 3174
rect 2384 3178 2444 4684
rect 3050 3722 3110 4684
rect 2854 3456 2930 3466
rect 2664 3450 2930 3456
rect 2740 3390 2762 3450
rect 2834 3390 2860 3450
rect 2928 3390 2930 3450
rect 2664 3384 2930 3390
rect 2854 3374 2930 3384
rect 1279 2166 1339 3118
rect 1718 2084 1776 3174
rect 1946 2084 2004 3174
rect 2384 2166 2444 3118
rect 2612 2084 2670 3174
rect 3050 2166 3110 3662
rect -364 2078 14 2084
rect -364 2018 -352 2078
rect -292 2018 -254 2078
rect -194 2018 -156 2078
rect -96 2018 -58 2078
rect 2 2018 14 2078
rect -364 2012 14 2018
rect 372 2078 1142 2084
rect 372 2018 384 2078
rect 444 2018 482 2078
rect 542 2018 580 2078
rect 640 2018 678 2078
rect 738 2018 776 2078
rect 836 2018 874 2078
rect 934 2018 972 2078
rect 1032 2018 1070 2078
rect 1130 2018 1142 2078
rect 372 2012 1142 2018
rect 1474 2078 2244 2084
rect 1474 2018 1486 2078
rect 1546 2018 1584 2078
rect 1644 2018 1682 2078
rect 1742 2018 1780 2078
rect 1840 2018 1878 2078
rect 1938 2018 1976 2078
rect 2036 2018 2074 2078
rect 2134 2018 2172 2078
rect 2232 2018 2244 2078
rect 1474 2012 2244 2018
rect 2612 2078 2892 2084
rect 2612 2018 2624 2078
rect 2684 2018 2722 2078
rect 2782 2018 2820 2078
rect 2880 2018 2892 2078
rect 2612 2012 2892 2018
<< viali >>
rect -352 4738 -292 4798
rect -254 4738 -194 4798
rect -156 4738 -96 4798
rect -58 4738 2 4798
rect 384 4738 444 4798
rect 482 4738 542 4798
rect 580 4738 640 4798
rect 678 4738 738 4798
rect 776 4738 836 4798
rect 874 4738 934 4798
rect 972 4738 1032 4798
rect 1070 4738 1130 4798
rect 1486 4738 1546 4798
rect 1584 4738 1644 4798
rect 1682 4738 1742 4798
rect 1780 4738 1840 4798
rect 1878 4738 1938 4798
rect 1976 4738 2036 4798
rect 2074 4738 2134 4798
rect 2172 4738 2232 4798
rect 2624 4738 2684 4798
rect 2722 4738 2782 4798
rect 2820 4738 2880 4798
rect 175 3662 235 3722
rect -210 3390 -194 3450
rect -194 3390 -150 3450
rect -112 3390 -100 3450
rect -100 3390 -52 3450
rect -14 3390 -6 3450
rect -6 3390 46 3450
rect 364 3390 416 3450
rect 416 3390 424 3450
rect 462 3390 510 3450
rect 510 3390 522 3450
rect 560 3390 604 3450
rect 604 3390 620 3450
rect 894 3390 910 3450
rect 910 3390 954 3450
rect 992 3390 1004 3450
rect 1004 3390 1052 3450
rect 1090 3390 1098 3450
rect 1098 3390 1150 3450
rect 1468 3390 1520 3450
rect 1520 3390 1528 3450
rect 1566 3390 1614 3450
rect 1614 3390 1626 3450
rect 1664 3390 1708 3450
rect 1708 3390 1724 3450
rect 1998 3390 2014 3450
rect 2014 3390 2058 3450
rect 2096 3390 2108 3450
rect 2108 3390 2156 3450
rect 2194 3390 2202 3450
rect 2202 3390 2254 3450
rect 1279 3118 1339 3178
rect 3050 3662 3110 3722
rect 2664 3390 2680 3450
rect 2680 3390 2724 3450
rect 2762 3390 2774 3450
rect 2774 3390 2822 3450
rect 2860 3390 2868 3450
rect 2868 3390 2920 3450
rect 2384 3118 2444 3178
rect -352 2018 -292 2078
rect -254 2018 -194 2078
rect -156 2018 -96 2078
rect -58 2018 2 2078
rect 384 2018 444 2078
rect 482 2018 542 2078
rect 580 2018 640 2078
rect 678 2018 738 2078
rect 776 2018 836 2078
rect 874 2018 934 2078
rect 972 2018 1032 2078
rect 1070 2018 1130 2078
rect 1486 2018 1546 2078
rect 1584 2018 1644 2078
rect 1682 2018 1742 2078
rect 1780 2018 1840 2078
rect 1878 2018 1938 2078
rect 1976 2018 2036 2078
rect 2074 2018 2134 2078
rect 2172 2018 2232 2078
rect 2624 2018 2684 2078
rect 2722 2018 2782 2078
rect 2820 2018 2880 2078
<< metal1 >>
rect -400 4798 3246 4816
rect -400 4738 -352 4798
rect -292 4738 -254 4798
rect -194 4738 -156 4798
rect -96 4738 -58 4798
rect 2 4738 384 4798
rect 444 4738 482 4798
rect 542 4738 580 4798
rect 640 4738 678 4798
rect 738 4738 776 4798
rect 836 4738 874 4798
rect 934 4738 972 4798
rect 1032 4738 1070 4798
rect 1130 4738 1486 4798
rect 1546 4738 1584 4798
rect 1644 4738 1682 4798
rect 1742 4738 1780 4798
rect 1840 4738 1878 4798
rect 1938 4738 1976 4798
rect 2036 4738 2074 4798
rect 2134 4738 2172 4798
rect 2232 4738 2624 4798
rect 2684 4738 2722 4798
rect 2782 4738 2820 4798
rect 2880 4738 3246 4798
rect -400 4720 3246 4738
rect -400 3656 -28 3728
rect 163 3722 3246 3728
rect 163 3662 175 3722
rect 235 3662 3050 3722
rect 3110 3662 3246 3722
rect 163 3656 3246 3662
rect -100 3456 -28 3656
rect 2096 3456 2168 3656
rect -222 3450 632 3456
rect -222 3390 -210 3450
rect -150 3390 -112 3450
rect -52 3390 -14 3450
rect 46 3390 364 3450
rect 424 3390 462 3450
rect 522 3390 560 3450
rect 620 3390 632 3450
rect -222 3384 632 3390
rect 882 3450 1736 3456
rect 882 3390 894 3450
rect 954 3390 992 3450
rect 1052 3390 1090 3450
rect 1150 3390 1468 3450
rect 1528 3390 1566 3450
rect 1626 3390 1664 3450
rect 1724 3390 1736 3450
rect 882 3384 1736 3390
rect 1986 3450 2286 3456
rect 1986 3390 1998 3450
rect 2058 3390 2096 3450
rect 2156 3390 2194 3450
rect 2254 3390 2286 3450
rect 1986 3384 2286 3390
rect 2652 3450 2952 3456
rect 2652 3390 2664 3450
rect 2724 3390 2762 3450
rect 2822 3390 2860 3450
rect 2920 3390 2952 3450
rect 2652 3384 2952 3390
rect 1005 3184 1077 3384
rect 2762 3184 2834 3384
rect -400 3112 1077 3184
rect 1267 3178 3246 3184
rect 1267 3118 1279 3178
rect 1339 3118 2384 3178
rect 2444 3118 3246 3178
rect 1267 3112 3246 3118
rect -400 2078 3246 2096
rect -400 2018 -352 2078
rect -292 2018 -254 2078
rect -194 2018 -156 2078
rect -96 2018 -58 2078
rect 2 2018 384 2078
rect 444 2018 482 2078
rect 542 2018 580 2078
rect 640 2018 678 2078
rect 738 2018 776 2078
rect 836 2018 874 2078
rect 934 2018 972 2078
rect 1032 2018 1070 2078
rect 1130 2018 1486 2078
rect 1546 2018 1584 2078
rect 1644 2018 1682 2078
rect 1742 2018 1780 2078
rect 1840 2018 1878 2078
rect 1938 2018 1976 2078
rect 2036 2018 2074 2078
rect 2134 2018 2172 2078
rect 2232 2018 2624 2078
rect 2684 2018 2722 2078
rect 2782 2018 2820 2078
rect 2880 2018 3246 2078
rect -400 2000 3246 2018
use nfet_12  nfet_12_0
timestamp 1623239895
transform 1 0 -262 0 1 2170
box -138 -210 1072 1210
use nfet_12  nfet_12_1
timestamp 1623239895
transform 1 0 842 0 1 2170
box -138 -210 1072 1210
use nfet_34  nfet_34_0
timestamp 1623055983
transform 1 0 2004 0 1 2170
box -196 -210 576 1210
use nfet_34  nfet_34_1
timestamp 1623055983
transform 1 0 2670 0 1 2170
box -196 -210 576 1210
use pfet_12  pfet_12_0
timestamp 1623147612
transform 1 0 -204 0 1 3679
box -196 -220 1014 1155
use pfet_12  pfet_12_1
timestamp 1623147612
transform 1 0 900 0 1 3679
box -196 -220 1014 1155
use pfet_34  pfet_34_0
timestamp 1623147637
transform 1 0 1808 0 1 3460
box 0 -2 772 1374
use pfet_34  pfet_34_1
timestamp 1623147637
transform 1 0 2474 0 1 3460
box 0 -2 772 1374
<< labels >>
flabel metal1 s 1260 4720 1356 4816 1 FreeSans 100 0 0 0 vccd
flabel metal1 s 1260 2000 1356 2096 1 FreeSans 100 0 0 0 v_crt
flabel metal1 s -200 3112 -128 3184 1 FreeSans 100 0 0 0 inn
flabel metal1 s -200 3656 -128 3728 1 FreeSans 100 0 0 0 inp
flabel metal1 s 2974 3656 3046 3728 1 FreeSans 100 0 0 0 outp
flabel metal1 s 2974 3112 3046 3184 1 FreeSans 100 0 0 0 outn
flabel pwell s -400 3308 -328 3380 1 FreeSans 100 0 0 0 vssd
<< end >>
