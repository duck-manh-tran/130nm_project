magic
tech sky130A
timestamp 1637172953
<< pwell >>
rect 0 0 600 610
<< nmos >>
rect 95 100 285 500
rect 315 100 505 500
<< ndiff >>
rect 65 489 95 500
rect 65 471 71 489
rect 89 471 95 489
rect 65 453 95 471
rect 65 435 71 453
rect 89 435 95 453
rect 65 417 95 435
rect 65 399 71 417
rect 89 399 95 417
rect 65 381 95 399
rect 65 363 71 381
rect 89 363 95 381
rect 65 345 95 363
rect 65 327 71 345
rect 89 327 95 345
rect 65 309 95 327
rect 65 291 71 309
rect 89 291 95 309
rect 65 273 95 291
rect 65 255 71 273
rect 89 255 95 273
rect 65 237 95 255
rect 65 219 71 237
rect 89 219 95 237
rect 65 201 95 219
rect 65 183 71 201
rect 89 183 95 201
rect 65 165 95 183
rect 65 147 71 165
rect 89 147 95 165
rect 65 129 95 147
rect 65 111 71 129
rect 89 111 95 129
rect 65 100 95 111
rect 285 489 315 500
rect 285 471 291 489
rect 309 471 315 489
rect 285 453 315 471
rect 285 435 291 453
rect 309 435 315 453
rect 285 417 315 435
rect 285 399 291 417
rect 309 399 315 417
rect 285 381 315 399
rect 285 363 291 381
rect 309 363 315 381
rect 285 345 315 363
rect 285 327 291 345
rect 309 327 315 345
rect 285 309 315 327
rect 285 291 291 309
rect 309 291 315 309
rect 285 273 315 291
rect 285 255 291 273
rect 309 255 315 273
rect 285 237 315 255
rect 285 219 291 237
rect 309 219 315 237
rect 285 201 315 219
rect 285 183 291 201
rect 309 183 315 201
rect 285 165 315 183
rect 285 147 291 165
rect 309 147 315 165
rect 285 129 315 147
rect 285 111 291 129
rect 309 111 315 129
rect 285 100 315 111
rect 505 489 535 500
rect 505 471 511 489
rect 529 471 535 489
rect 505 453 535 471
rect 505 435 511 453
rect 529 435 535 453
rect 505 417 535 435
rect 505 399 511 417
rect 529 399 535 417
rect 505 381 535 399
rect 505 363 511 381
rect 529 363 535 381
rect 505 345 535 363
rect 505 327 511 345
rect 529 327 535 345
rect 505 309 535 327
rect 505 291 511 309
rect 529 291 535 309
rect 505 273 535 291
rect 505 255 511 273
rect 529 255 535 273
rect 505 237 535 255
rect 505 219 511 237
rect 529 219 535 237
rect 505 201 535 219
rect 505 183 511 201
rect 529 183 535 201
rect 505 165 535 183
rect 505 147 511 165
rect 529 147 535 165
rect 505 129 535 147
rect 505 111 511 129
rect 529 111 535 129
rect 505 100 535 111
<< ndiffc >>
rect 71 471 89 489
rect 71 435 89 453
rect 71 399 89 417
rect 71 363 89 381
rect 71 327 89 345
rect 71 291 89 309
rect 71 255 89 273
rect 71 219 89 237
rect 71 183 89 201
rect 71 147 89 165
rect 71 111 89 129
rect 291 471 309 489
rect 291 435 309 453
rect 291 399 309 417
rect 291 363 309 381
rect 291 327 309 345
rect 291 291 309 309
rect 291 255 309 273
rect 291 219 309 237
rect 291 183 309 201
rect 291 147 309 165
rect 291 111 309 129
rect 511 471 529 489
rect 511 435 529 453
rect 511 399 529 417
rect 511 363 529 381
rect 511 327 529 345
rect 511 291 529 309
rect 511 255 529 273
rect 511 219 529 237
rect 511 183 529 201
rect 511 147 529 165
rect 511 111 529 129
<< poly >>
rect 95 500 285 550
rect 315 500 505 550
rect 95 87 285 100
rect 315 87 505 100
<< locali >>
rect 65 489 95 502
rect 65 471 71 489
rect 89 471 95 489
rect 65 453 95 471
rect 65 435 71 453
rect 89 435 95 453
rect 65 417 95 435
rect 65 399 71 417
rect 89 399 95 417
rect 65 381 95 399
rect 65 363 71 381
rect 89 363 95 381
rect 65 345 95 363
rect 65 327 71 345
rect 89 327 95 345
rect 65 309 95 327
rect 65 291 71 309
rect 89 291 95 309
rect 65 273 95 291
rect 65 255 71 273
rect 89 255 95 273
rect 65 237 95 255
rect 65 219 71 237
rect 89 219 95 237
rect 65 201 95 219
rect 65 183 71 201
rect 89 183 95 201
rect 65 165 95 183
rect 65 147 71 165
rect 89 147 95 165
rect 65 129 95 147
rect 65 111 71 129
rect 89 111 95 129
rect 65 98 95 111
rect 285 489 315 502
rect 285 471 291 489
rect 309 471 315 489
rect 285 453 315 471
rect 285 435 291 453
rect 309 435 315 453
rect 285 417 315 435
rect 285 399 291 417
rect 309 399 315 417
rect 285 381 315 399
rect 285 363 291 381
rect 309 363 315 381
rect 285 345 315 363
rect 285 327 291 345
rect 309 327 315 345
rect 285 309 315 327
rect 285 291 291 309
rect 309 291 315 309
rect 285 273 315 291
rect 285 255 291 273
rect 309 255 315 273
rect 285 237 315 255
rect 285 219 291 237
rect 309 219 315 237
rect 285 201 315 219
rect 285 183 291 201
rect 309 183 315 201
rect 285 165 315 183
rect 285 147 291 165
rect 309 147 315 165
rect 285 129 315 147
rect 285 111 291 129
rect 309 111 315 129
rect 285 98 315 111
rect 505 489 535 502
rect 505 471 511 489
rect 529 471 535 489
rect 505 453 535 471
rect 505 435 511 453
rect 529 435 535 453
rect 505 417 535 435
rect 505 399 511 417
rect 529 399 535 417
rect 505 381 535 399
rect 505 363 511 381
rect 529 363 535 381
rect 505 345 535 363
rect 505 327 511 345
rect 529 327 535 345
rect 505 309 535 327
rect 505 291 511 309
rect 529 291 535 309
rect 505 273 535 291
rect 505 255 511 273
rect 529 255 535 273
rect 505 237 535 255
rect 505 219 511 237
rect 529 219 535 237
rect 505 201 535 219
rect 505 183 511 201
rect 529 183 535 201
rect 505 165 535 183
rect 505 147 511 165
rect 529 147 535 165
rect 505 129 535 147
rect 505 111 511 129
rect 529 111 535 129
rect 505 98 535 111
<< end >>
