magic
tech sky130A
timestamp 1637141615
<< nwell >>
rect 0 0 400 1000
<< pmos >>
rect 105 100 295 900
<< pdiff >>
rect 75 887 105 900
rect 75 869 81 887
rect 99 869 105 887
rect 75 851 105 869
rect 75 833 81 851
rect 99 833 105 851
rect 75 815 105 833
rect 75 797 81 815
rect 99 797 105 815
rect 75 779 105 797
rect 75 761 81 779
rect 99 761 105 779
rect 75 743 105 761
rect 75 725 81 743
rect 99 725 105 743
rect 75 707 105 725
rect 75 689 81 707
rect 99 689 105 707
rect 75 671 105 689
rect 75 653 81 671
rect 99 653 105 671
rect 75 635 105 653
rect 75 617 81 635
rect 99 617 105 635
rect 75 599 105 617
rect 75 581 81 599
rect 99 581 105 599
rect 75 563 105 581
rect 75 545 81 563
rect 99 545 105 563
rect 75 527 105 545
rect 75 509 81 527
rect 99 509 105 527
rect 75 491 105 509
rect 75 473 81 491
rect 99 473 105 491
rect 75 455 105 473
rect 75 437 81 455
rect 99 437 105 455
rect 75 419 105 437
rect 75 401 81 419
rect 99 401 105 419
rect 75 383 105 401
rect 75 365 81 383
rect 99 365 105 383
rect 75 347 105 365
rect 75 329 81 347
rect 99 329 105 347
rect 75 311 105 329
rect 75 293 81 311
rect 99 293 105 311
rect 75 275 105 293
rect 75 257 81 275
rect 99 257 105 275
rect 75 239 105 257
rect 75 221 81 239
rect 99 221 105 239
rect 75 203 105 221
rect 75 185 81 203
rect 99 185 105 203
rect 75 167 105 185
rect 75 149 81 167
rect 99 149 105 167
rect 75 131 105 149
rect 75 113 81 131
rect 99 113 105 131
rect 75 100 105 113
rect 295 887 325 900
rect 295 869 301 887
rect 319 869 325 887
rect 295 851 325 869
rect 295 833 301 851
rect 319 833 325 851
rect 295 815 325 833
rect 295 797 301 815
rect 319 797 325 815
rect 295 779 325 797
rect 295 761 301 779
rect 319 761 325 779
rect 295 743 325 761
rect 295 725 301 743
rect 319 725 325 743
rect 295 707 325 725
rect 295 689 301 707
rect 319 689 325 707
rect 295 671 325 689
rect 295 653 301 671
rect 319 653 325 671
rect 295 635 325 653
rect 295 617 301 635
rect 319 617 325 635
rect 295 599 325 617
rect 295 581 301 599
rect 319 581 325 599
rect 295 563 325 581
rect 295 545 301 563
rect 319 545 325 563
rect 295 527 325 545
rect 295 509 301 527
rect 319 509 325 527
rect 295 491 325 509
rect 295 473 301 491
rect 319 473 325 491
rect 295 455 325 473
rect 295 437 301 455
rect 319 437 325 455
rect 295 419 325 437
rect 295 401 301 419
rect 319 401 325 419
rect 295 383 325 401
rect 295 365 301 383
rect 319 365 325 383
rect 295 347 325 365
rect 295 329 301 347
rect 319 329 325 347
rect 295 311 325 329
rect 295 293 301 311
rect 319 293 325 311
rect 295 275 325 293
rect 295 257 301 275
rect 319 257 325 275
rect 295 239 325 257
rect 295 221 301 239
rect 319 221 325 239
rect 295 203 325 221
rect 295 185 301 203
rect 319 185 325 203
rect 295 167 325 185
rect 295 149 301 167
rect 319 149 325 167
rect 295 131 325 149
rect 295 113 301 131
rect 319 113 325 131
rect 295 100 325 113
<< pdiffc >>
rect 81 869 99 887
rect 81 833 99 851
rect 81 797 99 815
rect 81 761 99 779
rect 81 725 99 743
rect 81 689 99 707
rect 81 653 99 671
rect 81 617 99 635
rect 81 581 99 599
rect 81 545 99 563
rect 81 509 99 527
rect 81 473 99 491
rect 81 437 99 455
rect 81 401 99 419
rect 81 365 99 383
rect 81 329 99 347
rect 81 293 99 311
rect 81 257 99 275
rect 81 221 99 239
rect 81 185 99 203
rect 81 149 99 167
rect 81 113 99 131
rect 301 869 319 887
rect 301 833 319 851
rect 301 797 319 815
rect 301 761 319 779
rect 301 725 319 743
rect 301 689 319 707
rect 301 653 319 671
rect 301 617 319 635
rect 301 581 319 599
rect 301 545 319 563
rect 301 509 319 527
rect 301 473 319 491
rect 301 437 319 455
rect 301 401 319 419
rect 301 365 319 383
rect 301 329 319 347
rect 301 293 319 311
rect 301 257 319 275
rect 301 221 319 239
rect 301 185 319 203
rect 301 149 319 167
rect 301 113 319 131
<< nsubdiff >>
rect 35 934 47 952
rect 65 934 83 952
rect 101 934 119 952
rect 137 934 155 952
rect 173 934 191 952
rect 209 934 227 952
rect 245 934 263 952
rect 281 934 299 952
rect 317 934 335 952
rect 353 934 365 952
<< nsubdiffcont >>
rect 47 934 65 952
rect 83 934 101 952
rect 119 934 137 952
rect 155 934 173 952
rect 191 934 209 952
rect 227 934 245 952
rect 263 934 281 952
rect 299 934 317 952
rect 335 934 353 952
<< poly >>
rect 105 900 295 913
rect 105 52 295 100
<< locali >>
rect 35 934 47 952
rect 65 934 83 952
rect 101 934 119 952
rect 137 934 155 952
rect 173 934 191 952
rect 209 934 227 952
rect 245 934 263 952
rect 281 934 299 952
rect 317 934 335 952
rect 353 934 365 952
rect 75 887 105 934
rect 75 869 81 887
rect 99 869 105 887
rect 75 851 105 869
rect 75 833 81 851
rect 99 833 105 851
rect 75 815 105 833
rect 75 797 81 815
rect 99 797 105 815
rect 75 779 105 797
rect 75 761 81 779
rect 99 761 105 779
rect 75 743 105 761
rect 75 725 81 743
rect 99 725 105 743
rect 75 707 105 725
rect 75 689 81 707
rect 99 689 105 707
rect 75 671 105 689
rect 75 653 81 671
rect 99 653 105 671
rect 75 635 105 653
rect 75 617 81 635
rect 99 617 105 635
rect 75 599 105 617
rect 75 581 81 599
rect 99 581 105 599
rect 75 563 105 581
rect 75 545 81 563
rect 99 545 105 563
rect 75 527 105 545
rect 75 509 81 527
rect 99 509 105 527
rect 75 491 105 509
rect 75 473 81 491
rect 99 473 105 491
rect 75 455 105 473
rect 75 437 81 455
rect 99 437 105 455
rect 75 419 105 437
rect 75 401 81 419
rect 99 401 105 419
rect 75 383 105 401
rect 75 365 81 383
rect 99 365 105 383
rect 75 347 105 365
rect 75 329 81 347
rect 99 329 105 347
rect 75 311 105 329
rect 75 293 81 311
rect 99 293 105 311
rect 75 275 105 293
rect 75 257 81 275
rect 99 257 105 275
rect 75 239 105 257
rect 75 221 81 239
rect 99 221 105 239
rect 75 203 105 221
rect 75 185 81 203
rect 99 185 105 203
rect 75 167 105 185
rect 75 149 81 167
rect 99 149 105 167
rect 75 131 105 149
rect 75 113 81 131
rect 99 113 105 131
rect 75 98 105 113
rect 295 887 325 902
rect 295 869 301 887
rect 319 869 325 887
rect 295 851 325 869
rect 295 833 301 851
rect 319 833 325 851
rect 295 815 325 833
rect 295 797 301 815
rect 319 797 325 815
rect 295 779 325 797
rect 295 761 301 779
rect 319 761 325 779
rect 295 743 325 761
rect 295 725 301 743
rect 319 725 325 743
rect 295 707 325 725
rect 295 689 301 707
rect 319 689 325 707
rect 295 671 325 689
rect 295 653 301 671
rect 319 653 325 671
rect 295 635 325 653
rect 295 617 301 635
rect 319 617 325 635
rect 295 599 325 617
rect 295 581 301 599
rect 319 581 325 599
rect 295 563 325 581
rect 295 545 301 563
rect 319 545 325 563
rect 295 527 325 545
rect 295 509 301 527
rect 319 509 325 527
rect 295 491 325 509
rect 295 473 301 491
rect 319 473 325 491
rect 295 455 325 473
rect 295 437 301 455
rect 319 437 325 455
rect 295 419 325 437
rect 295 401 301 419
rect 319 401 325 419
rect 295 383 325 401
rect 295 365 301 383
rect 319 365 325 383
rect 295 347 325 365
rect 295 329 301 347
rect 319 329 325 347
rect 295 311 325 329
rect 295 293 301 311
rect 319 293 325 311
rect 295 275 325 293
rect 295 257 301 275
rect 319 257 325 275
rect 295 239 325 257
rect 295 221 301 239
rect 319 221 325 239
rect 295 203 325 221
rect 295 185 301 203
rect 319 185 325 203
rect 295 167 325 185
rect 295 149 301 167
rect 319 149 325 167
rect 295 131 325 149
rect 295 113 301 131
rect 319 113 325 131
rect 295 98 325 113
<< end >>
