magic
tech sky130A
timestamp 1637401559
<< poly >>
rect 69 636 479 684
rect 69 619 75 636
rect 92 619 111 636
rect 128 619 147 636
rect 164 619 183 636
rect 200 619 348 636
rect 365 619 384 636
rect 401 619 420 636
rect 437 619 456 636
rect 473 619 479 636
rect 69 599 479 619
rect 69 582 75 599
rect 92 582 111 599
rect 128 582 147 599
rect 164 582 183 599
rect 200 582 348 599
rect 365 582 384 599
rect 401 582 420 599
rect 437 582 456 599
rect 473 582 479 599
rect 69 534 479 582
rect 617 636 1027 684
rect 617 619 623 636
rect 640 619 659 636
rect 676 619 695 636
rect 712 619 731 636
rect 748 619 896 636
rect 913 619 932 636
rect 949 619 968 636
rect 985 619 1004 636
rect 1021 619 1027 636
rect 617 599 1027 619
rect 617 582 623 599
rect 640 582 659 599
rect 676 582 695 599
rect 712 582 731 599
rect 748 582 896 599
rect 913 582 932 599
rect 949 582 968 599
rect 985 582 1004 599
rect 1021 582 1027 599
rect 617 534 1027 582
rect 1165 636 1355 686
rect 1165 619 1171 636
rect 1188 619 1207 636
rect 1224 619 1243 636
rect 1260 619 1279 636
rect 1296 619 1355 636
rect 1165 599 1355 619
rect 1165 582 1171 599
rect 1188 582 1207 599
rect 1224 582 1243 599
rect 1260 582 1279 599
rect 1296 582 1355 599
rect 1165 528 1355 582
rect 1453 636 1643 686
rect 1453 619 1459 636
rect 1476 619 1495 636
rect 1512 619 1531 636
rect 1548 619 1567 636
rect 1584 619 1643 636
rect 1453 599 1643 619
rect 1453 582 1459 599
rect 1476 582 1495 599
rect 1512 582 1531 599
rect 1548 582 1567 599
rect 1584 582 1643 599
rect 1453 528 1643 582
<< polycont >>
rect 75 619 92 636
rect 111 619 128 636
rect 147 619 164 636
rect 183 619 200 636
rect 348 619 365 636
rect 384 619 401 636
rect 420 619 437 636
rect 456 619 473 636
rect 75 582 92 599
rect 111 582 128 599
rect 147 582 164 599
rect 183 582 200 599
rect 348 582 365 599
rect 384 582 401 599
rect 420 582 437 599
rect 456 582 473 599
rect 623 619 640 636
rect 659 619 676 636
rect 695 619 712 636
rect 731 619 748 636
rect 896 619 913 636
rect 932 619 949 636
rect 968 619 985 636
rect 1004 619 1021 636
rect 623 582 640 599
rect 659 582 676 599
rect 695 582 712 599
rect 731 582 748 599
rect 896 582 913 599
rect 932 582 949 599
rect 968 582 985 599
rect 1004 582 1021 599
rect 1171 619 1188 636
rect 1207 619 1224 636
rect 1243 619 1260 636
rect 1279 619 1296 636
rect 1171 582 1188 599
rect 1207 582 1224 599
rect 1243 582 1260 599
rect 1279 582 1296 599
rect 1459 619 1476 636
rect 1495 619 1512 636
rect 1531 619 1548 636
rect 1567 619 1584 636
rect 1459 582 1476 599
rect 1495 582 1512 599
rect 1531 582 1548 599
rect 1567 582 1584 599
<< locali >>
rect -9 1581 11 1605
rect 35 1581 82 1605
rect 106 1581 154 1605
rect 178 1581 226 1605
rect 250 1581 298 1605
rect 322 1581 370 1605
rect 394 1581 442 1605
rect 466 1581 514 1605
rect 538 1581 594 1605
rect 618 1581 666 1605
rect 690 1581 738 1605
rect 762 1581 810 1605
rect 834 1581 882 1605
rect 906 1581 954 1605
rect 978 1581 1026 1605
rect 1050 1581 1104 1605
rect 1128 1581 1176 1605
rect 1200 1581 1248 1605
rect 1272 1581 1320 1605
rect 1344 1581 1392 1605
rect 1416 1581 1464 1605
rect 1488 1581 1536 1605
rect 1560 1581 1608 1605
rect 1632 1581 1679 1605
rect 1703 1581 1712 1605
rect 259 749 289 769
rect 259 731 265 749
rect 283 731 289 749
rect 67 619 75 636
rect 92 619 111 636
rect 128 619 147 636
rect 164 619 183 636
rect 200 619 208 636
rect 67 582 75 599
rect 92 582 111 599
rect 128 582 147 599
rect 164 582 183 599
rect 200 582 208 599
rect 259 480 289 731
rect 340 619 348 636
rect 365 619 384 636
rect 401 619 420 636
rect 437 619 456 636
rect 473 619 481 636
rect 615 619 623 636
rect 640 619 659 636
rect 676 619 695 636
rect 712 619 731 636
rect 748 619 756 636
rect 340 582 348 599
rect 365 582 384 599
rect 401 582 420 599
rect 437 582 456 599
rect 473 582 481 599
rect 615 582 623 599
rect 640 582 659 599
rect 676 582 695 599
rect 712 582 731 599
rect 748 582 756 599
rect 807 487 837 733
rect 888 619 896 636
rect 913 619 932 636
rect 949 619 968 636
rect 985 619 1004 636
rect 1021 619 1029 636
rect 1163 619 1171 636
rect 1188 619 1207 636
rect 1224 619 1243 636
rect 1260 619 1279 636
rect 1296 619 1304 636
rect 888 582 896 599
rect 913 582 932 599
rect 949 582 968 599
rect 985 582 1004 599
rect 1021 582 1029 599
rect 1163 582 1171 599
rect 1188 582 1207 599
rect 1224 582 1243 599
rect 1260 582 1279 599
rect 1296 582 1304 599
rect 807 469 813 487
rect 831 469 837 487
rect 1355 486 1385 777
rect 1643 769 1649 786
rect 1667 769 1673 786
rect 1643 749 1673 769
rect 1643 731 1649 749
rect 1667 731 1673 749
rect 1451 619 1459 636
rect 1476 619 1495 636
rect 1512 619 1531 636
rect 1548 619 1567 636
rect 1584 619 1592 636
rect 1451 582 1459 599
rect 1476 582 1495 599
rect 1512 582 1531 599
rect 1548 582 1567 599
rect 1584 582 1592 599
rect 1355 468 1361 486
rect 1379 468 1385 486
rect 1355 449 1385 468
rect 807 432 813 449
rect 831 432 837 449
rect 1355 432 1361 449
rect 1379 432 1385 449
rect 1643 435 1673 731
rect 39 38 69 82
rect 479 38 509 82
rect 587 38 617 82
rect 1027 38 1057 82
rect 1135 38 1165 82
rect 1423 38 1453 82
rect 0 12 10 38
rect 36 12 66 38
rect 92 12 122 38
rect 148 12 178 38
rect 204 12 234 38
rect 260 12 290 38
rect 316 12 346 38
rect 372 12 402 38
rect 428 12 458 38
rect 484 12 514 38
rect 540 12 570 38
rect 596 12 626 38
rect 652 12 682 38
rect 708 12 738 38
rect 764 12 794 38
rect 820 12 850 38
rect 876 12 906 38
rect 932 12 962 38
rect 988 12 1018 38
rect 1044 12 1074 38
rect 1100 12 1130 38
rect 1156 12 1186 38
rect 1212 12 1242 38
rect 1268 12 1298 38
rect 1324 12 1354 38
rect 1380 12 1410 38
rect 1436 12 1466 38
rect 1492 12 1522 38
rect 1548 12 1578 38
rect 1604 12 1634 38
rect 1660 12 1712 38
<< viali >>
rect 11 1581 35 1605
rect 82 1581 106 1605
rect 154 1581 178 1605
rect 226 1581 250 1605
rect 298 1581 322 1605
rect 370 1581 394 1605
rect 442 1581 466 1605
rect 514 1581 538 1605
rect 594 1581 618 1605
rect 666 1581 690 1605
rect 738 1581 762 1605
rect 810 1581 834 1605
rect 882 1581 906 1605
rect 954 1581 978 1605
rect 1026 1581 1050 1605
rect 1104 1581 1128 1605
rect 1176 1581 1200 1605
rect 1248 1581 1272 1605
rect 1320 1581 1344 1605
rect 1392 1581 1416 1605
rect 1464 1581 1488 1605
rect 1536 1581 1560 1605
rect 1608 1581 1632 1605
rect 1679 1581 1703 1605
rect 265 769 283 787
rect 265 731 283 749
rect 75 619 92 636
rect 111 619 128 636
rect 147 619 164 636
rect 183 619 200 636
rect 75 582 92 599
rect 111 582 128 599
rect 147 582 164 599
rect 183 582 200 599
rect 348 619 365 636
rect 384 619 401 636
rect 420 619 437 636
rect 456 619 473 636
rect 623 619 640 636
rect 659 619 676 636
rect 695 619 712 636
rect 731 619 748 636
rect 348 582 365 599
rect 384 582 401 599
rect 420 582 437 599
rect 456 582 473 599
rect 623 582 640 599
rect 659 582 676 599
rect 695 582 712 599
rect 731 582 748 599
rect 896 619 913 636
rect 932 619 949 636
rect 968 619 985 636
rect 1004 619 1021 636
rect 1171 619 1188 636
rect 1207 619 1224 636
rect 1243 619 1260 636
rect 1279 619 1296 636
rect 896 582 913 599
rect 932 582 949 599
rect 968 582 985 599
rect 1004 582 1021 599
rect 1171 582 1188 599
rect 1207 582 1224 599
rect 1243 582 1260 599
rect 1279 582 1296 599
rect 813 469 831 487
rect 1649 769 1667 787
rect 1649 731 1667 749
rect 1459 619 1476 636
rect 1495 619 1512 636
rect 1531 619 1548 636
rect 1567 619 1584 636
rect 1459 582 1476 599
rect 1495 582 1512 599
rect 1531 582 1548 599
rect 1567 582 1584 599
rect 1361 468 1379 486
rect 813 431 831 449
rect 1361 431 1379 449
rect 10 12 36 38
rect 66 12 92 38
rect 122 12 148 38
rect 178 12 204 38
rect 234 12 260 38
rect 290 12 316 38
rect 346 12 372 38
rect 402 12 428 38
rect 458 12 484 38
rect 514 12 540 38
rect 570 12 596 38
rect 626 12 652 38
rect 682 12 708 38
rect 738 12 764 38
rect 794 12 820 38
rect 850 12 876 38
rect 906 12 932 38
rect 962 12 988 38
rect 1018 12 1044 38
rect 1074 12 1100 38
rect 1130 12 1156 38
rect 1186 12 1212 38
rect 1242 12 1268 38
rect 1298 12 1324 38
rect 1354 12 1380 38
rect 1410 12 1436 38
rect 1466 12 1492 38
rect 1522 12 1548 38
rect 1578 12 1604 38
rect 1634 12 1660 38
<< metal1 >>
rect -9 1605 1712 1619
rect -9 1581 11 1605
rect 35 1581 82 1605
rect 106 1581 154 1605
rect 178 1581 226 1605
rect 250 1581 298 1605
rect 322 1581 370 1605
rect 394 1581 442 1605
rect 466 1581 514 1605
rect 538 1581 594 1605
rect 618 1581 666 1605
rect 690 1581 738 1605
rect 762 1581 810 1605
rect 834 1581 882 1605
rect 906 1581 954 1605
rect 978 1581 1026 1605
rect 1050 1581 1104 1605
rect 1128 1581 1176 1605
rect 1200 1581 1248 1605
rect 1272 1581 1320 1605
rect 1344 1581 1392 1605
rect 1416 1581 1464 1605
rect 1488 1581 1536 1605
rect 1560 1581 1608 1605
rect 1632 1581 1679 1605
rect 1703 1581 1712 1605
rect -9 1569 1712 1581
rect 259 787 289 790
rect 0 734 174 784
rect 124 639 174 734
rect 259 769 265 787
rect 283 784 289 787
rect 1643 787 1673 790
rect 1643 784 1649 787
rect 283 769 1649 784
rect 1667 784 1673 787
rect 1667 769 1712 784
rect 259 749 1712 769
rect 259 731 265 749
rect 283 734 1649 749
rect 283 731 289 734
rect 259 728 289 731
rect 1224 639 1274 734
rect 1643 731 1649 734
rect 1667 734 1712 749
rect 1667 731 1673 734
rect 1643 728 1673 731
rect 69 636 208 639
rect 69 619 75 636
rect 92 619 111 636
rect 128 619 147 636
rect 164 619 183 636
rect 200 634 208 636
rect 340 636 479 639
rect 340 634 348 636
rect 200 619 348 634
rect 365 619 384 636
rect 401 619 420 636
rect 437 619 456 636
rect 473 619 479 636
rect 69 599 479 619
rect 69 582 75 599
rect 92 582 111 599
rect 128 582 147 599
rect 164 582 183 599
rect 200 584 348 599
rect 200 582 208 584
rect 69 579 208 582
rect 340 582 348 584
rect 365 582 384 599
rect 401 582 420 599
rect 437 582 456 599
rect 473 582 479 599
rect 340 579 479 582
rect 617 636 756 639
rect 617 619 623 636
rect 640 619 659 636
rect 676 619 695 636
rect 712 619 731 636
rect 748 634 756 636
rect 888 636 1027 639
rect 888 634 896 636
rect 748 619 896 634
rect 913 619 932 636
rect 949 619 968 636
rect 985 619 1004 636
rect 1021 619 1027 636
rect 617 599 1027 619
rect 617 582 623 599
rect 640 582 659 599
rect 676 582 695 599
rect 712 582 731 599
rect 748 584 896 599
rect 748 582 756 584
rect 617 579 756 582
rect 888 582 896 584
rect 913 582 932 599
rect 949 582 968 599
rect 985 582 1004 599
rect 1021 582 1027 599
rect 888 579 1027 582
rect 1165 636 1304 639
rect 1165 619 1171 636
rect 1188 619 1207 636
rect 1224 619 1243 636
rect 1260 619 1279 636
rect 1296 619 1304 636
rect 1165 599 1304 619
rect 1165 582 1171 599
rect 1188 582 1207 599
rect 1224 582 1243 599
rect 1260 582 1279 599
rect 1296 582 1304 599
rect 1165 579 1304 582
rect 1453 636 1592 639
rect 1453 619 1459 636
rect 1476 619 1495 636
rect 1512 619 1531 636
rect 1548 619 1567 636
rect 1584 619 1592 636
rect 1453 599 1592 619
rect 1453 582 1459 599
rect 1476 582 1495 599
rect 1512 582 1531 599
rect 1548 582 1567 599
rect 1584 582 1592 599
rect 1453 579 1592 582
rect 674 484 724 579
rect 0 434 724 484
rect 807 487 837 490
rect 807 469 813 487
rect 831 484 837 487
rect 1355 486 1385 490
rect 1355 484 1361 486
rect 831 469 1361 484
rect 807 468 1361 469
rect 1379 484 1385 486
rect 1508 484 1558 579
rect 1379 468 1712 484
rect 807 449 1712 468
rect 807 431 813 449
rect 831 434 1361 449
rect 831 431 837 434
rect 807 428 837 431
rect 1355 431 1361 434
rect 1379 434 1712 449
rect 1379 431 1385 434
rect 1355 428 1385 431
rect 0 38 1712 50
rect 0 12 10 38
rect 36 12 66 38
rect 92 12 122 38
rect 148 12 178 38
rect 204 12 234 38
rect 260 12 290 38
rect 316 12 346 38
rect 372 12 402 38
rect 428 12 458 38
rect 484 12 514 38
rect 540 12 570 38
rect 596 12 626 38
rect 652 12 682 38
rect 708 12 738 38
rect 764 12 794 38
rect 820 12 850 38
rect 876 12 906 38
rect 932 12 962 38
rect 988 12 1018 38
rect 1044 12 1074 38
rect 1100 12 1130 38
rect 1156 12 1186 38
rect 1212 12 1242 38
rect 1268 12 1298 38
rect 1324 12 1354 38
rect 1380 12 1410 38
rect 1436 12 1466 38
rect 1492 12 1522 38
rect 1548 12 1578 38
rect 1604 12 1634 38
rect 1660 12 1712 38
rect 0 0 1712 12
use nfet_12  nfet_12_0
timestamp 1637401559
transform 1 0 -26 0 1 -16
box 0 0 600 610
use nfet_12  nfet_12_1
timestamp 1637401559
transform 1 0 522 0 1 -16
box 0 0 600 610
use pfet_12  pfet_12_0
timestamp 1637401559
transform 1 0 -76 0 1 634
box 0 0 700 1016
use nfet_34  nfet_34_0
timestamp 1637401559
transform 1 0 1060 0 1 -16
box 0 0 400 610
use nfet_34  nfet_34_1
timestamp 1637401559
transform 1 0 1348 0 1 -16
box 0 0 400 610
use pfet_34  pfet_34_0
timestamp 1637401559
transform 1 0 1060 0 1 634
box 0 0 400 1016
use pfet_34  pfet_34_1
timestamp 1637401559
transform 1 0 1348 0 1 634
box 0 0 400 1016
use pfet_12  pfet_12_1
timestamp 1637401559
transform 1 0 472 0 1 634
box 0 0 700 1016
<< labels >>
flabel metal1 16 760 16 760 1 FreeSans 240 0 0 0 inn
flabel metal1 18 459 18 459 1 FreeSans 240 0 0 0 inp
flabel metal1 1100 760 1100 760 1 FreeSans 240 0 0 0 outn
flabel metal1 1100 459 1100 459 1 FreeSans 240 0 0 0 outp
<< end >>
