magic
tech sky130A
timestamp 1623170494
<< metal3 >>
rect 15300 12780 29900 12800
rect 15300 12740 15320 12780
rect 15360 12740 15380 12780
rect 15420 12740 15440 12780
rect 15480 12740 18920 12780
rect 18960 12740 18980 12780
rect 19020 12740 19040 12780
rect 19080 12740 22520 12780
rect 22560 12740 22580 12780
rect 22620 12740 22640 12780
rect 22680 12740 26120 12780
rect 26160 12740 26180 12780
rect 26220 12740 26240 12780
rect 26280 12740 29720 12780
rect 29760 12740 29780 12780
rect 29820 12740 29840 12780
rect 29880 12740 29900 12780
rect 15300 12720 29900 12740
rect 15300 12680 15320 12720
rect 15360 12680 15380 12720
rect 15420 12680 15440 12720
rect 15480 12680 18920 12720
rect 18960 12680 18980 12720
rect 19020 12680 19040 12720
rect 19080 12680 22520 12720
rect 22560 12680 22580 12720
rect 22620 12680 22640 12720
rect 22680 12680 26120 12720
rect 26160 12680 26180 12720
rect 26220 12680 26240 12720
rect 26280 12680 29720 12720
rect 29760 12680 29780 12720
rect 29820 12680 29840 12720
rect 29880 12680 29900 12720
rect 15300 12660 29900 12680
rect 15300 12620 15320 12660
rect 15360 12620 15380 12660
rect 15420 12620 15440 12660
rect 15480 12620 18920 12660
rect 18960 12620 18980 12660
rect 19020 12620 19040 12660
rect 19080 12620 22520 12660
rect 22560 12620 22580 12660
rect 22620 12620 22640 12660
rect 22680 12620 26120 12660
rect 26160 12620 26180 12660
rect 26220 12620 26240 12660
rect 26280 12620 29720 12660
rect 29760 12620 29780 12660
rect 29820 12620 29840 12660
rect 29880 12620 29900 12660
rect 15300 12600 29900 12620
rect 13500 12180 31700 12200
rect 13500 12140 13520 12180
rect 13560 12140 13580 12180
rect 13620 12140 13640 12180
rect 13680 12140 17120 12180
rect 17160 12140 17180 12180
rect 17220 12140 17240 12180
rect 17280 12140 20720 12180
rect 20760 12140 20780 12180
rect 20820 12140 20840 12180
rect 20880 12140 24320 12180
rect 24360 12140 24380 12180
rect 24420 12140 24440 12180
rect 24480 12140 27920 12180
rect 27960 12140 27980 12180
rect 28020 12140 28040 12180
rect 28080 12140 31520 12180
rect 31560 12140 31580 12180
rect 31620 12140 31640 12180
rect 31680 12140 31700 12180
rect 13500 12120 31700 12140
rect 13500 12080 13520 12120
rect 13560 12080 13580 12120
rect 13620 12080 13640 12120
rect 13680 12080 17120 12120
rect 17160 12080 17180 12120
rect 17220 12080 17240 12120
rect 17280 12080 20720 12120
rect 20760 12080 20780 12120
rect 20820 12080 20840 12120
rect 20880 12080 24320 12120
rect 24360 12080 24380 12120
rect 24420 12080 24440 12120
rect 24480 12080 27920 12120
rect 27960 12080 27980 12120
rect 28020 12080 28040 12120
rect 28080 12080 31520 12120
rect 31560 12080 31580 12120
rect 31620 12080 31640 12120
rect 31680 12080 31700 12120
rect 13500 12060 31700 12080
rect 13500 12020 13520 12060
rect 13560 12020 13580 12060
rect 13620 12020 13640 12060
rect 13680 12020 17120 12060
rect 17160 12020 17180 12060
rect 17220 12020 17240 12060
rect 17280 12020 20720 12060
rect 20760 12020 20780 12060
rect 20820 12020 20840 12060
rect 20880 12020 24320 12060
rect 24360 12020 24380 12060
rect 24420 12020 24440 12060
rect 24480 12020 27920 12060
rect 27960 12020 27980 12060
rect 28020 12020 28040 12060
rect 28080 12020 31520 12060
rect 31560 12020 31580 12060
rect 31620 12020 31640 12060
rect 31680 12020 31700 12060
rect 13500 12000 31700 12020
rect 13500 1680 31700 1700
rect 13500 1640 13520 1680
rect 13560 1640 13580 1680
rect 13620 1640 13640 1680
rect 13680 1640 17120 1680
rect 17160 1640 17180 1680
rect 17220 1640 17240 1680
rect 17280 1640 20720 1680
rect 20760 1640 20780 1680
rect 20820 1640 20840 1680
rect 20880 1640 24320 1680
rect 24360 1640 24380 1680
rect 24420 1640 24440 1680
rect 24480 1640 27920 1680
rect 27960 1640 27980 1680
rect 28020 1640 28040 1680
rect 28080 1640 31520 1680
rect 31560 1640 31580 1680
rect 31620 1640 31640 1680
rect 31680 1640 31700 1680
rect 13500 1620 31700 1640
rect 13500 1580 13520 1620
rect 13560 1580 13580 1620
rect 13620 1580 13640 1620
rect 13680 1580 17120 1620
rect 17160 1580 17180 1620
rect 17220 1580 17240 1620
rect 17280 1580 20720 1620
rect 20760 1580 20780 1620
rect 20820 1580 20840 1620
rect 20880 1580 24320 1620
rect 24360 1580 24380 1620
rect 24420 1580 24440 1620
rect 24480 1580 27920 1620
rect 27960 1580 27980 1620
rect 28020 1580 28040 1620
rect 28080 1580 31520 1620
rect 31560 1580 31580 1620
rect 31620 1580 31640 1620
rect 31680 1580 31700 1620
rect 13500 1560 31700 1580
rect 13500 1520 13520 1560
rect 13560 1520 13580 1560
rect 13620 1520 13640 1560
rect 13680 1520 17120 1560
rect 17160 1520 17180 1560
rect 17220 1520 17240 1560
rect 17280 1520 20720 1560
rect 20760 1520 20780 1560
rect 20820 1520 20840 1560
rect 20880 1520 24320 1560
rect 24360 1520 24380 1560
rect 24420 1520 24440 1560
rect 24480 1520 27920 1560
rect 27960 1520 27980 1560
rect 28020 1520 28040 1560
rect 28080 1520 31520 1560
rect 31560 1520 31580 1560
rect 31620 1520 31640 1560
rect 31680 1520 31700 1560
rect 13500 1500 31700 1520
rect 15300 1080 29900 1100
rect 15300 1040 15320 1080
rect 15360 1040 15380 1080
rect 15420 1040 15440 1080
rect 15480 1040 18920 1080
rect 18960 1040 18980 1080
rect 19020 1040 19040 1080
rect 19080 1040 22520 1080
rect 22560 1040 22580 1080
rect 22620 1040 22640 1080
rect 22680 1040 26120 1080
rect 26160 1040 26180 1080
rect 26220 1040 26240 1080
rect 26280 1040 29720 1080
rect 29760 1040 29780 1080
rect 29820 1040 29840 1080
rect 29880 1040 29900 1080
rect 15300 1020 29900 1040
rect 15300 980 15320 1020
rect 15360 980 15380 1020
rect 15420 980 15440 1020
rect 15480 980 18920 1020
rect 18960 980 18980 1020
rect 19020 980 19040 1020
rect 19080 980 22520 1020
rect 22560 980 22580 1020
rect 22620 980 22640 1020
rect 22680 980 26120 1020
rect 26160 980 26180 1020
rect 26220 980 26240 1020
rect 26280 980 29720 1020
rect 29760 980 29780 1020
rect 29820 980 29840 1020
rect 29880 980 29900 1020
rect 15300 960 29900 980
rect 15300 920 15320 960
rect 15360 920 15380 960
rect 15420 920 15440 960
rect 15480 920 18920 960
rect 18960 920 18980 960
rect 19020 920 19040 960
rect 19080 920 22520 960
rect 22560 920 22580 960
rect 22620 920 22640 960
rect 22680 920 26120 960
rect 26160 920 26180 960
rect 26220 920 26240 960
rect 26280 920 29720 960
rect 29760 920 29780 960
rect 29820 920 29840 960
rect 29880 920 29900 960
rect 15300 900 29900 920
<< via3 >>
rect 15320 12740 15360 12780
rect 15380 12740 15420 12780
rect 15440 12740 15480 12780
rect 18920 12740 18960 12780
rect 18980 12740 19020 12780
rect 19040 12740 19080 12780
rect 22520 12740 22560 12780
rect 22580 12740 22620 12780
rect 22640 12740 22680 12780
rect 26120 12740 26160 12780
rect 26180 12740 26220 12780
rect 26240 12740 26280 12780
rect 29720 12740 29760 12780
rect 29780 12740 29820 12780
rect 29840 12740 29880 12780
rect 15320 12680 15360 12720
rect 15380 12680 15420 12720
rect 15440 12680 15480 12720
rect 18920 12680 18960 12720
rect 18980 12680 19020 12720
rect 19040 12680 19080 12720
rect 22520 12680 22560 12720
rect 22580 12680 22620 12720
rect 22640 12680 22680 12720
rect 26120 12680 26160 12720
rect 26180 12680 26220 12720
rect 26240 12680 26280 12720
rect 29720 12680 29760 12720
rect 29780 12680 29820 12720
rect 29840 12680 29880 12720
rect 15320 12620 15360 12660
rect 15380 12620 15420 12660
rect 15440 12620 15480 12660
rect 18920 12620 18960 12660
rect 18980 12620 19020 12660
rect 19040 12620 19080 12660
rect 22520 12620 22560 12660
rect 22580 12620 22620 12660
rect 22640 12620 22680 12660
rect 26120 12620 26160 12660
rect 26180 12620 26220 12660
rect 26240 12620 26280 12660
rect 29720 12620 29760 12660
rect 29780 12620 29820 12660
rect 29840 12620 29880 12660
rect 13520 12140 13560 12180
rect 13580 12140 13620 12180
rect 13640 12140 13680 12180
rect 17120 12140 17160 12180
rect 17180 12140 17220 12180
rect 17240 12140 17280 12180
rect 20720 12140 20760 12180
rect 20780 12140 20820 12180
rect 20840 12140 20880 12180
rect 24320 12140 24360 12180
rect 24380 12140 24420 12180
rect 24440 12140 24480 12180
rect 27920 12140 27960 12180
rect 27980 12140 28020 12180
rect 28040 12140 28080 12180
rect 31520 12140 31560 12180
rect 31580 12140 31620 12180
rect 31640 12140 31680 12180
rect 13520 12080 13560 12120
rect 13580 12080 13620 12120
rect 13640 12080 13680 12120
rect 17120 12080 17160 12120
rect 17180 12080 17220 12120
rect 17240 12080 17280 12120
rect 20720 12080 20760 12120
rect 20780 12080 20820 12120
rect 20840 12080 20880 12120
rect 24320 12080 24360 12120
rect 24380 12080 24420 12120
rect 24440 12080 24480 12120
rect 27920 12080 27960 12120
rect 27980 12080 28020 12120
rect 28040 12080 28080 12120
rect 31520 12080 31560 12120
rect 31580 12080 31620 12120
rect 31640 12080 31680 12120
rect 13520 12020 13560 12060
rect 13580 12020 13620 12060
rect 13640 12020 13680 12060
rect 17120 12020 17160 12060
rect 17180 12020 17220 12060
rect 17240 12020 17280 12060
rect 20720 12020 20760 12060
rect 20780 12020 20820 12060
rect 20840 12020 20880 12060
rect 24320 12020 24360 12060
rect 24380 12020 24420 12060
rect 24440 12020 24480 12060
rect 27920 12020 27960 12060
rect 27980 12020 28020 12060
rect 28040 12020 28080 12060
rect 31520 12020 31560 12060
rect 31580 12020 31620 12060
rect 31640 12020 31680 12060
rect 13520 1640 13560 1680
rect 13580 1640 13620 1680
rect 13640 1640 13680 1680
rect 17120 1640 17160 1680
rect 17180 1640 17220 1680
rect 17240 1640 17280 1680
rect 20720 1640 20760 1680
rect 20780 1640 20820 1680
rect 20840 1640 20880 1680
rect 24320 1640 24360 1680
rect 24380 1640 24420 1680
rect 24440 1640 24480 1680
rect 27920 1640 27960 1680
rect 27980 1640 28020 1680
rect 28040 1640 28080 1680
rect 31520 1640 31560 1680
rect 31580 1640 31620 1680
rect 31640 1640 31680 1680
rect 13520 1580 13560 1620
rect 13580 1580 13620 1620
rect 13640 1580 13680 1620
rect 17120 1580 17160 1620
rect 17180 1580 17220 1620
rect 17240 1580 17280 1620
rect 20720 1580 20760 1620
rect 20780 1580 20820 1620
rect 20840 1580 20880 1620
rect 24320 1580 24360 1620
rect 24380 1580 24420 1620
rect 24440 1580 24480 1620
rect 27920 1580 27960 1620
rect 27980 1580 28020 1620
rect 28040 1580 28080 1620
rect 31520 1580 31560 1620
rect 31580 1580 31620 1620
rect 31640 1580 31680 1620
rect 13520 1520 13560 1560
rect 13580 1520 13620 1560
rect 13640 1520 13680 1560
rect 17120 1520 17160 1560
rect 17180 1520 17220 1560
rect 17240 1520 17280 1560
rect 20720 1520 20760 1560
rect 20780 1520 20820 1560
rect 20840 1520 20880 1560
rect 24320 1520 24360 1560
rect 24380 1520 24420 1560
rect 24440 1520 24480 1560
rect 27920 1520 27960 1560
rect 27980 1520 28020 1560
rect 28040 1520 28080 1560
rect 31520 1520 31560 1560
rect 31580 1520 31620 1560
rect 31640 1520 31680 1560
rect 15320 1040 15360 1080
rect 15380 1040 15420 1080
rect 15440 1040 15480 1080
rect 18920 1040 18960 1080
rect 18980 1040 19020 1080
rect 19040 1040 19080 1080
rect 22520 1040 22560 1080
rect 22580 1040 22620 1080
rect 22640 1040 22680 1080
rect 26120 1040 26160 1080
rect 26180 1040 26220 1080
rect 26240 1040 26280 1080
rect 29720 1040 29760 1080
rect 29780 1040 29820 1080
rect 29840 1040 29880 1080
rect 15320 980 15360 1020
rect 15380 980 15420 1020
rect 15440 980 15480 1020
rect 18920 980 18960 1020
rect 18980 980 19020 1020
rect 19040 980 19080 1020
rect 22520 980 22560 1020
rect 22580 980 22620 1020
rect 22640 980 22680 1020
rect 26120 980 26160 1020
rect 26180 980 26220 1020
rect 26240 980 26280 1020
rect 29720 980 29760 1020
rect 29780 980 29820 1020
rect 29840 980 29880 1020
rect 15320 920 15360 960
rect 15380 920 15420 960
rect 15440 920 15480 960
rect 18920 920 18960 960
rect 18980 920 19020 960
rect 19040 920 19080 960
rect 22520 920 22560 960
rect 22580 920 22620 960
rect 22640 920 22680 960
rect 26120 920 26160 960
rect 26180 920 26220 960
rect 26240 920 26280 960
rect 29720 920 29760 960
rect 29780 920 29820 960
rect 29840 920 29880 960
<< metal4 >>
rect 15300 12780 15500 12800
rect 15300 12740 15320 12780
rect 15360 12740 15380 12780
rect 15420 12740 15440 12780
rect 15480 12740 15500 12780
rect 15300 12720 15500 12740
rect 15300 12680 15320 12720
rect 15360 12680 15380 12720
rect 15420 12680 15440 12720
rect 15480 12680 15500 12720
rect 15300 12660 15500 12680
rect 15300 12620 15320 12660
rect 15360 12620 15380 12660
rect 15420 12620 15440 12660
rect 15480 12620 15500 12660
rect 13500 12180 13700 12200
rect 13500 12140 13520 12180
rect 13560 12140 13580 12180
rect 13620 12140 13640 12180
rect 13680 12140 13700 12180
rect 13500 12120 13700 12140
rect 13500 12080 13520 12120
rect 13560 12080 13580 12120
rect 13620 12080 13640 12120
rect 13680 12080 13700 12120
rect 13500 12060 13700 12080
rect 13500 12020 13520 12060
rect 13560 12020 13580 12060
rect 13620 12020 13640 12060
rect 13680 12020 13700 12060
rect 13500 1680 13700 12020
rect 13500 1640 13520 1680
rect 13560 1640 13580 1680
rect 13620 1640 13640 1680
rect 13680 1640 13700 1680
rect 13500 1620 13700 1640
rect 13500 1580 13520 1620
rect 13560 1580 13580 1620
rect 13620 1580 13640 1620
rect 13680 1580 13700 1620
rect 13500 1560 13700 1580
rect 13500 1520 13520 1560
rect 13560 1520 13580 1560
rect 13620 1520 13640 1560
rect 13680 1520 13700 1560
rect 13500 1500 13700 1520
rect 15300 1080 15500 12620
rect 18900 12780 19100 12800
rect 18900 12740 18920 12780
rect 18960 12740 18980 12780
rect 19020 12740 19040 12780
rect 19080 12740 19100 12780
rect 18900 12720 19100 12740
rect 18900 12680 18920 12720
rect 18960 12680 18980 12720
rect 19020 12680 19040 12720
rect 19080 12680 19100 12720
rect 18900 12660 19100 12680
rect 18900 12620 18920 12660
rect 18960 12620 18980 12660
rect 19020 12620 19040 12660
rect 19080 12620 19100 12660
rect 17100 12180 17300 12200
rect 17100 12140 17120 12180
rect 17160 12140 17180 12180
rect 17220 12140 17240 12180
rect 17280 12140 17300 12180
rect 17100 12120 17300 12140
rect 17100 12080 17120 12120
rect 17160 12080 17180 12120
rect 17220 12080 17240 12120
rect 17280 12080 17300 12120
rect 17100 12060 17300 12080
rect 17100 12020 17120 12060
rect 17160 12020 17180 12060
rect 17220 12020 17240 12060
rect 17280 12020 17300 12060
rect 17100 8900 17300 12020
rect 17100 1680 17300 4750
rect 17100 1640 17120 1680
rect 17160 1640 17180 1680
rect 17220 1640 17240 1680
rect 17280 1640 17300 1680
rect 17100 1620 17300 1640
rect 17100 1580 17120 1620
rect 17160 1580 17180 1620
rect 17220 1580 17240 1620
rect 17280 1580 17300 1620
rect 17100 1560 17300 1580
rect 17100 1520 17120 1560
rect 17160 1520 17180 1560
rect 17220 1520 17240 1560
rect 17280 1520 17300 1560
rect 17100 1500 17300 1520
rect 15300 1040 15320 1080
rect 15360 1040 15380 1080
rect 15420 1040 15440 1080
rect 15480 1040 15500 1080
rect 15300 1020 15500 1040
rect 15300 980 15320 1020
rect 15360 980 15380 1020
rect 15420 980 15440 1020
rect 15480 980 15500 1020
rect 15300 960 15500 980
rect 15300 920 15320 960
rect 15360 920 15380 960
rect 15420 920 15440 960
rect 15480 920 15500 960
rect 15300 900 15500 920
rect 18900 1080 19100 12620
rect 22500 12780 22700 12800
rect 22500 12740 22520 12780
rect 22560 12740 22580 12780
rect 22620 12740 22640 12780
rect 22680 12740 22700 12780
rect 22500 12720 22700 12740
rect 22500 12680 22520 12720
rect 22560 12680 22580 12720
rect 22620 12680 22640 12720
rect 22680 12680 22700 12720
rect 22500 12660 22700 12680
rect 22500 12620 22520 12660
rect 22560 12620 22580 12660
rect 22620 12620 22640 12660
rect 22680 12620 22700 12660
rect 20700 12180 20900 12200
rect 20700 12140 20720 12180
rect 20760 12140 20780 12180
rect 20820 12140 20840 12180
rect 20880 12140 20900 12180
rect 20700 12120 20900 12140
rect 20700 12080 20720 12120
rect 20760 12080 20780 12120
rect 20820 12080 20840 12120
rect 20880 12080 20900 12120
rect 20700 12060 20900 12080
rect 20700 12020 20720 12060
rect 20760 12020 20780 12060
rect 20820 12020 20840 12060
rect 20880 12020 20900 12060
rect 20700 8900 20900 12020
rect 20700 1680 20900 4750
rect 20700 1640 20720 1680
rect 20760 1640 20780 1680
rect 20820 1640 20840 1680
rect 20880 1640 20900 1680
rect 20700 1620 20900 1640
rect 20700 1580 20720 1620
rect 20760 1580 20780 1620
rect 20820 1580 20840 1620
rect 20880 1580 20900 1620
rect 20700 1560 20900 1580
rect 20700 1520 20720 1560
rect 20760 1520 20780 1560
rect 20820 1520 20840 1560
rect 20880 1520 20900 1560
rect 20700 1500 20900 1520
rect 18900 1040 18920 1080
rect 18960 1040 18980 1080
rect 19020 1040 19040 1080
rect 19080 1040 19100 1080
rect 18900 1020 19100 1040
rect 18900 980 18920 1020
rect 18960 980 18980 1020
rect 19020 980 19040 1020
rect 19080 980 19100 1020
rect 18900 960 19100 980
rect 18900 920 18920 960
rect 18960 920 18980 960
rect 19020 920 19040 960
rect 19080 920 19100 960
rect 18900 900 19100 920
rect 22500 1080 22700 12620
rect 26100 12780 26300 12800
rect 26100 12740 26120 12780
rect 26160 12740 26180 12780
rect 26220 12740 26240 12780
rect 26280 12740 26300 12780
rect 26100 12720 26300 12740
rect 26100 12680 26120 12720
rect 26160 12680 26180 12720
rect 26220 12680 26240 12720
rect 26280 12680 26300 12720
rect 26100 12660 26300 12680
rect 26100 12620 26120 12660
rect 26160 12620 26180 12660
rect 26220 12620 26240 12660
rect 26280 12620 26300 12660
rect 24300 12180 24500 12200
rect 24300 12140 24320 12180
rect 24360 12140 24380 12180
rect 24420 12140 24440 12180
rect 24480 12140 24500 12180
rect 24300 12120 24500 12140
rect 24300 12080 24320 12120
rect 24360 12080 24380 12120
rect 24420 12080 24440 12120
rect 24480 12080 24500 12120
rect 24300 12060 24500 12080
rect 24300 12020 24320 12060
rect 24360 12020 24380 12060
rect 24420 12020 24440 12060
rect 24480 12020 24500 12060
rect 24300 8900 24500 12020
rect 24300 1680 24500 4750
rect 24300 1640 24320 1680
rect 24360 1640 24380 1680
rect 24420 1640 24440 1680
rect 24480 1640 24500 1680
rect 24300 1620 24500 1640
rect 24300 1580 24320 1620
rect 24360 1580 24380 1620
rect 24420 1580 24440 1620
rect 24480 1580 24500 1620
rect 24300 1560 24500 1580
rect 24300 1520 24320 1560
rect 24360 1520 24380 1560
rect 24420 1520 24440 1560
rect 24480 1520 24500 1560
rect 24300 1500 24500 1520
rect 22500 1040 22520 1080
rect 22560 1040 22580 1080
rect 22620 1040 22640 1080
rect 22680 1040 22700 1080
rect 22500 1020 22700 1040
rect 22500 980 22520 1020
rect 22560 980 22580 1020
rect 22620 980 22640 1020
rect 22680 980 22700 1020
rect 22500 960 22700 980
rect 22500 920 22520 960
rect 22560 920 22580 960
rect 22620 920 22640 960
rect 22680 920 22700 960
rect 22500 900 22700 920
rect 26100 1080 26300 12620
rect 29700 12780 29900 12800
rect 29700 12740 29720 12780
rect 29760 12740 29780 12780
rect 29820 12740 29840 12780
rect 29880 12740 29900 12780
rect 29700 12720 29900 12740
rect 29700 12680 29720 12720
rect 29760 12680 29780 12720
rect 29820 12680 29840 12720
rect 29880 12680 29900 12720
rect 29700 12660 29900 12680
rect 29700 12620 29720 12660
rect 29760 12620 29780 12660
rect 29820 12620 29840 12660
rect 29880 12620 29900 12660
rect 27900 12180 28100 12200
rect 27900 12140 27920 12180
rect 27960 12140 27980 12180
rect 28020 12140 28040 12180
rect 28080 12140 28100 12180
rect 27900 12120 28100 12140
rect 27900 12080 27920 12120
rect 27960 12080 27980 12120
rect 28020 12080 28040 12120
rect 28080 12080 28100 12120
rect 27900 12060 28100 12080
rect 27900 12020 27920 12060
rect 27960 12020 27980 12060
rect 28020 12020 28040 12060
rect 28080 12020 28100 12060
rect 27900 8900 28100 12020
rect 27900 1680 28100 4750
rect 27900 1640 27920 1680
rect 27960 1640 27980 1680
rect 28020 1640 28040 1680
rect 28080 1640 28100 1680
rect 27900 1620 28100 1640
rect 27900 1580 27920 1620
rect 27960 1580 27980 1620
rect 28020 1580 28040 1620
rect 28080 1580 28100 1620
rect 27900 1560 28100 1580
rect 27900 1520 27920 1560
rect 27960 1520 27980 1560
rect 28020 1520 28040 1560
rect 28080 1520 28100 1560
rect 27900 1500 28100 1520
rect 26100 1040 26120 1080
rect 26160 1040 26180 1080
rect 26220 1040 26240 1080
rect 26280 1040 26300 1080
rect 26100 1020 26300 1040
rect 26100 980 26120 1020
rect 26160 980 26180 1020
rect 26220 980 26240 1020
rect 26280 980 26300 1020
rect 26100 960 26300 980
rect 26100 920 26120 960
rect 26160 920 26180 960
rect 26220 920 26240 960
rect 26280 920 26300 960
rect 26100 900 26300 920
rect 29700 1080 29900 12620
rect 31500 12180 31700 12200
rect 31500 12140 31520 12180
rect 31560 12140 31580 12180
rect 31620 12140 31640 12180
rect 31680 12140 31700 12180
rect 31500 12120 31700 12140
rect 31500 12080 31520 12120
rect 31560 12080 31580 12120
rect 31620 12080 31640 12120
rect 31680 12080 31700 12120
rect 31500 12060 31700 12080
rect 31500 12020 31520 12060
rect 31560 12020 31580 12060
rect 31620 12020 31640 12060
rect 31680 12020 31700 12060
rect 31500 1680 31700 12020
rect 31500 1640 31520 1680
rect 31560 1640 31580 1680
rect 31620 1640 31640 1680
rect 31680 1640 31700 1680
rect 31500 1620 31700 1640
rect 31500 1580 31520 1620
rect 31560 1580 31580 1620
rect 31620 1580 31640 1620
rect 31680 1580 31700 1620
rect 31500 1560 31700 1580
rect 31500 1520 31520 1560
rect 31560 1520 31580 1560
rect 31620 1520 31640 1560
rect 31680 1520 31700 1560
rect 31500 1500 31700 1520
rect 29700 1040 29720 1080
rect 29760 1040 29780 1080
rect 29820 1040 29840 1080
rect 29880 1040 29900 1080
rect 29700 1020 29900 1040
rect 29700 980 29720 1020
rect 29760 980 29780 1020
rect 29820 980 29840 1020
rect 29880 980 29900 1020
rect 29700 960 29900 980
rect 29700 920 29720 960
rect 29760 920 29780 960
rect 29820 920 29840 960
rect 29880 920 29900 960
rect 29700 900 29900 920
<< end >>
