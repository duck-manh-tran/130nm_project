magic
tech sky130A
magscale 1 2
timestamp 1623644919
<< nwell >>
rect -200 5142 336 5190
rect -162 5120 38 5142
<< nsubdiff >>
rect -162 5120 -122 5154
rect -82 5120 -42 5154
rect -2 5120 38 5154
<< nsubdiffcont >>
rect -122 5120 -82 5154
rect -42 5120 -2 5154
<< poly >>
rect 20500 3900 20600 3973
rect 20500 3878 20673 3900
rect 20500 3832 20532 3878
rect 20578 3832 20673 3878
rect 20500 3800 20673 3832
<< polycont >>
rect 20532 3832 20578 3878
<< locali >>
rect -162 5120 -122 5154
rect -82 5120 -42 5154
rect -2 5120 38 5154
rect 336 4950 601 4992
rect 281 4948 601 4950
rect 281 4906 380 4948
rect 557 4907 601 4948
rect 557 4863 654 4907
rect 442 4856 502 4862
rect 442 4808 448 4856
rect 496 4808 502 4856
rect 442 4696 502 4808
rect 281 4636 502 4696
rect 20400 3900 20600 3973
rect 20400 3884 20673 3900
rect 20400 3824 20418 3884
rect 20478 3824 20522 3884
rect 20582 3824 20673 3884
rect 20400 3780 20673 3824
rect 20400 3720 20418 3780
rect 20478 3720 20522 3780
rect 20582 3720 20673 3780
rect 20400 3700 20673 3720
rect 21504 3880 21700 3900
rect 21504 3875 21521 3880
rect 21504 3820 21519 3875
rect 21581 3820 21619 3880
rect 21679 3820 21700 3880
rect 21504 3780 21700 3820
rect 21504 3720 21521 3780
rect 21581 3720 21619 3780
rect 21679 3720 21700 3780
rect 21504 3700 21700 3720
<< viali >>
rect 448 4808 496 4856
rect 20220 4810 20280 4870
rect 20320 4810 20380 4870
rect 20420 4810 20480 4870
rect 20520 4810 20580 4870
rect 20418 3824 20478 3884
rect 20522 3878 20582 3884
rect 20522 3832 20532 3878
rect 20532 3832 20578 3878
rect 20578 3832 20582 3878
rect 20522 3824 20582 3832
rect 20418 3720 20478 3780
rect 20522 3720 20582 3780
rect 21521 3820 21581 3880
rect 21619 3820 21679 3880
rect 21521 3720 21581 3780
rect 21619 3720 21679 3780
<< metal1 >>
rect 1680 5854 1914 5950
rect -200 5056 640 5152
rect 20200 4870 20601 4876
rect 436 4856 1698 4862
rect 436 4808 448 4856
rect 496 4808 1698 4856
rect 436 4802 1698 4808
rect 1152 4790 1698 4802
rect 5254 4790 5326 4862
rect 8796 4790 8868 4862
rect 12334 4790 12406 4862
rect 15878 4790 15950 4862
rect 19508 4790 20044 4862
rect 20200 4810 20220 4870
rect 20280 4810 20320 4870
rect 20380 4810 20420 4870
rect 20480 4810 20520 4870
rect 20580 4810 20601 4870
rect 20200 4803 20601 4810
rect -200 4512 637 4608
rect 1152 3472 1224 4790
rect -502 3400 1224 3472
rect 1424 4246 1702 4318
rect 5254 4246 5326 4318
rect 8798 4246 8870 4318
rect 12334 4246 12406 4318
rect 15878 4246 15950 4318
rect 19504 4246 19772 4318
rect -502 1178 -430 3400
rect 1424 3200 1496 4246
rect -230 3128 1496 3200
rect 2400 3206 2600 3230
rect 2452 3154 2474 3206
rect 2526 3154 2548 3206
rect 2400 3134 2600 3154
rect 3600 3206 3800 3230
rect 3652 3154 3674 3206
rect 3726 3154 3748 3206
rect 3600 3134 3800 3154
rect 4800 3206 5000 3230
rect 4852 3154 4874 3206
rect 4926 3154 4948 3206
rect 4800 3134 5000 3154
rect 6000 3206 6200 3230
rect 6052 3154 6074 3206
rect 6126 3154 6148 3206
rect 6000 3134 6200 3154
rect 7200 3206 7400 3230
rect 7252 3154 7274 3206
rect 7326 3154 7348 3206
rect 7200 3134 7400 3154
rect 8400 3206 8600 3230
rect 8452 3154 8474 3206
rect 8526 3154 8548 3206
rect 8400 3134 8600 3154
rect 9600 3206 9800 3230
rect 9652 3154 9674 3206
rect 9726 3154 9748 3206
rect 9600 3134 9800 3154
rect 10800 3206 11000 3230
rect 10852 3154 10874 3206
rect 10926 3154 10948 3206
rect 10800 3134 11000 3154
rect 12000 3206 12200 3230
rect 12052 3154 12074 3206
rect 12126 3154 12148 3206
rect 12000 3134 12200 3154
rect 13200 3206 13400 3230
rect 13252 3154 13274 3206
rect 13326 3154 13348 3206
rect 13200 3134 13400 3154
rect 14400 3206 14600 3230
rect 14452 3154 14474 3206
rect 14526 3154 14548 3206
rect 14400 3134 14600 3154
rect 15600 3206 15800 3230
rect 15652 3154 15674 3206
rect 15726 3154 15748 3206
rect 15600 3134 15800 3154
rect 16800 3206 17000 3230
rect 16852 3154 16874 3206
rect 16926 3154 16948 3206
rect 16800 3134 17000 3154
rect 18000 3206 18200 3230
rect 18052 3154 18074 3206
rect 18126 3154 18148 3206
rect 18000 3134 18200 3154
rect 19200 3206 19400 3230
rect 19252 3154 19274 3206
rect 19326 3154 19348 3206
rect 19200 3134 19400 3154
rect 19700 3200 19772 4246
rect 19972 3472 20044 4790
rect 20400 3888 20600 3903
rect 20400 3820 20414 3888
rect 20482 3820 20518 3888
rect 20586 3820 20600 3888
rect 20400 3784 20600 3820
rect 20400 3716 20414 3784
rect 20482 3716 20518 3784
rect 20586 3716 20600 3784
rect 20400 3700 20600 3716
rect 21503 3884 21700 3900
rect 21503 3816 21517 3884
rect 21585 3816 21615 3884
rect 21683 3816 21700 3884
rect 21503 3784 21700 3816
rect 21503 3716 21517 3784
rect 21585 3716 21615 3784
rect 21683 3716 21700 3784
rect 21503 3700 21700 3716
rect 19972 3400 21872 3472
rect 19700 3128 21600 3200
rect -230 1722 -158 3128
rect 0 2810 200 2834
rect 52 2758 74 2810
rect 126 2758 148 2810
rect 0 2738 200 2758
rect 1200 2810 1400 2834
rect 1252 2758 1274 2810
rect 1326 2758 1348 2810
rect 1200 2738 1400 2758
rect 2400 2810 2600 2834
rect 2452 2758 2474 2810
rect 2526 2758 2548 2810
rect 2400 2738 2600 2758
rect 3600 2810 3800 2834
rect 3652 2758 3674 2810
rect 3726 2758 3748 2810
rect 3600 2738 3800 2758
rect 4800 2810 5000 2834
rect 4852 2758 4874 2810
rect 4926 2758 4948 2810
rect 4800 2738 5000 2758
rect 6000 2810 6200 2834
rect 6052 2758 6074 2810
rect 6126 2758 6148 2810
rect 6000 2738 6200 2758
rect 7200 2810 7400 2834
rect 7252 2758 7274 2810
rect 7326 2758 7348 2810
rect 7200 2738 7400 2758
rect 8400 2810 8600 2834
rect 8452 2758 8474 2810
rect 8526 2758 8548 2810
rect 8400 2738 8600 2758
rect 9600 2810 9800 2834
rect 9652 2758 9674 2810
rect 9726 2758 9748 2810
rect 9600 2738 9800 2758
rect 10800 2810 11000 2834
rect 10852 2758 10874 2810
rect 10926 2758 10948 2810
rect 10800 2738 11000 2758
rect 12000 2810 12200 2834
rect 12052 2758 12074 2810
rect 12126 2758 12148 2810
rect 12000 2738 12200 2758
rect 13200 2810 13400 2834
rect 13252 2758 13274 2810
rect 13326 2758 13348 2810
rect 13200 2738 13400 2758
rect 14400 2810 14600 2834
rect 14452 2758 14474 2810
rect 14526 2758 14548 2810
rect 14400 2738 14600 2758
rect 15600 2810 15800 2834
rect 15652 2758 15674 2810
rect 15726 2758 15748 2810
rect 15600 2738 15800 2758
rect 16800 2810 17000 2834
rect 16852 2758 16874 2810
rect 16926 2758 16948 2810
rect 16800 2738 17000 2758
rect 18000 2810 18200 2834
rect 18052 2758 18074 2810
rect 18126 2758 18148 2810
rect 18000 2738 18200 2758
rect 19200 2810 19400 2834
rect 19252 2758 19274 2810
rect 19326 2758 19348 2810
rect 19200 2738 19400 2758
rect 20400 2810 20600 2834
rect 20452 2758 20474 2810
rect 20526 2758 20548 2810
rect 20400 2738 20600 2758
rect 21156 2810 21356 2834
rect 21208 2758 21230 2810
rect 21282 2758 21304 2810
rect 21156 2738 21356 2758
rect 21528 1722 21600 3128
rect -230 1650 0 1722
rect 3554 1650 3626 1722
rect 7104 1650 7176 1722
rect 10634 1650 10706 1722
rect 14182 1650 14254 1722
rect 17728 1650 17800 1722
rect 21267 1650 21600 1722
rect 21800 1178 21872 3400
rect -502 1106 0 1178
rect 3556 1106 3628 1178
rect 7106 1106 7178 1178
rect 10650 1106 10722 1178
rect 14182 1106 14254 1178
rect 17728 1106 17802 1178
rect 21356 1106 21872 1178
<< via1 >>
rect 2400 3154 2452 3206
rect 2474 3154 2526 3206
rect 2548 3154 2600 3206
rect 3600 3154 3652 3206
rect 3674 3154 3726 3206
rect 3748 3154 3800 3206
rect 4800 3154 4852 3206
rect 4874 3154 4926 3206
rect 4948 3154 5000 3206
rect 6000 3154 6052 3206
rect 6074 3154 6126 3206
rect 6148 3154 6200 3206
rect 7200 3154 7252 3206
rect 7274 3154 7326 3206
rect 7348 3154 7400 3206
rect 8400 3154 8452 3206
rect 8474 3154 8526 3206
rect 8548 3154 8600 3206
rect 9600 3154 9652 3206
rect 9674 3154 9726 3206
rect 9748 3154 9800 3206
rect 10800 3154 10852 3206
rect 10874 3154 10926 3206
rect 10948 3154 11000 3206
rect 12000 3154 12052 3206
rect 12074 3154 12126 3206
rect 12148 3154 12200 3206
rect 13200 3154 13252 3206
rect 13274 3154 13326 3206
rect 13348 3154 13400 3206
rect 14400 3154 14452 3206
rect 14474 3154 14526 3206
rect 14548 3154 14600 3206
rect 15600 3154 15652 3206
rect 15674 3154 15726 3206
rect 15748 3154 15800 3206
rect 16800 3154 16852 3206
rect 16874 3154 16926 3206
rect 16948 3154 17000 3206
rect 18000 3154 18052 3206
rect 18074 3154 18126 3206
rect 18148 3154 18200 3206
rect 19200 3154 19252 3206
rect 19274 3154 19326 3206
rect 19348 3154 19400 3206
rect 20414 3884 20482 3888
rect 20414 3824 20418 3884
rect 20418 3824 20478 3884
rect 20478 3824 20482 3884
rect 20414 3820 20482 3824
rect 20518 3884 20586 3888
rect 20518 3824 20522 3884
rect 20522 3824 20582 3884
rect 20582 3824 20586 3884
rect 20518 3820 20586 3824
rect 20414 3780 20482 3784
rect 20414 3720 20418 3780
rect 20418 3720 20478 3780
rect 20478 3720 20482 3780
rect 20414 3716 20482 3720
rect 20518 3780 20586 3784
rect 20518 3720 20522 3780
rect 20522 3720 20582 3780
rect 20582 3720 20586 3780
rect 20518 3716 20586 3720
rect 21517 3880 21585 3884
rect 21517 3820 21521 3880
rect 21521 3820 21581 3880
rect 21581 3820 21585 3880
rect 21517 3816 21585 3820
rect 21615 3880 21683 3884
rect 21615 3820 21619 3880
rect 21619 3820 21679 3880
rect 21679 3820 21683 3880
rect 21615 3816 21683 3820
rect 21517 3780 21585 3784
rect 21517 3720 21521 3780
rect 21521 3720 21581 3780
rect 21581 3720 21585 3780
rect 21517 3716 21585 3720
rect 21615 3780 21683 3784
rect 21615 3720 21619 3780
rect 21619 3720 21679 3780
rect 21679 3720 21683 3780
rect 21615 3716 21683 3720
rect 0 2758 52 2810
rect 74 2758 126 2810
rect 148 2758 200 2810
rect 1200 2758 1252 2810
rect 1274 2758 1326 2810
rect 1348 2758 1400 2810
rect 2400 2758 2452 2810
rect 2474 2758 2526 2810
rect 2548 2758 2600 2810
rect 3600 2758 3652 2810
rect 3674 2758 3726 2810
rect 3748 2758 3800 2810
rect 4800 2758 4852 2810
rect 4874 2758 4926 2810
rect 4948 2758 5000 2810
rect 6000 2758 6052 2810
rect 6074 2758 6126 2810
rect 6148 2758 6200 2810
rect 7200 2758 7252 2810
rect 7274 2758 7326 2810
rect 7348 2758 7400 2810
rect 8400 2758 8452 2810
rect 8474 2758 8526 2810
rect 8548 2758 8600 2810
rect 9600 2758 9652 2810
rect 9674 2758 9726 2810
rect 9748 2758 9800 2810
rect 10800 2758 10852 2810
rect 10874 2758 10926 2810
rect 10948 2758 11000 2810
rect 12000 2758 12052 2810
rect 12074 2758 12126 2810
rect 12148 2758 12200 2810
rect 13200 2758 13252 2810
rect 13274 2758 13326 2810
rect 13348 2758 13400 2810
rect 14400 2758 14452 2810
rect 14474 2758 14526 2810
rect 14548 2758 14600 2810
rect 15600 2758 15652 2810
rect 15674 2758 15726 2810
rect 15748 2758 15800 2810
rect 16800 2758 16852 2810
rect 16874 2758 16926 2810
rect 16948 2758 17000 2810
rect 18000 2758 18052 2810
rect 18074 2758 18126 2810
rect 18148 2758 18200 2810
rect 19200 2758 19252 2810
rect 19274 2758 19326 2810
rect 19348 2758 19400 2810
rect 20400 2758 20452 2810
rect 20474 2758 20526 2810
rect 20548 2758 20600 2810
rect 21156 2758 21208 2810
rect 21230 2758 21282 2810
rect 21304 2758 21356 2810
<< metal2 >>
rect 20400 3894 20600 3903
rect 20400 3814 20408 3894
rect 20488 3814 20512 3894
rect 20592 3814 20600 3894
rect 20400 3790 20600 3814
rect 20400 3710 20408 3790
rect 20488 3710 20512 3790
rect 20592 3710 20600 3790
rect 20400 3700 20600 3710
rect 21503 3884 21700 3900
rect 21503 3816 21517 3884
rect 21585 3816 21615 3884
rect 21683 3816 21700 3884
rect 21503 3784 21700 3816
rect 21503 3716 21517 3784
rect 21585 3716 21615 3784
rect 21683 3716 21700 3784
rect 21503 3700 21700 3716
rect 2400 3210 2600 3220
rect 2400 3206 2420 3210
rect 2480 3206 2520 3210
rect 2580 3206 2600 3210
rect 2400 3150 2420 3154
rect 2480 3150 2520 3154
rect 2580 3150 2600 3154
rect 2400 3140 2600 3150
rect 3600 3210 3800 3220
rect 3600 3206 3620 3210
rect 3680 3206 3720 3210
rect 3780 3206 3800 3210
rect 3600 3150 3620 3154
rect 3680 3150 3720 3154
rect 3780 3150 3800 3154
rect 3600 3140 3800 3150
rect 4800 3210 5000 3220
rect 4800 3206 4820 3210
rect 4880 3206 4920 3210
rect 4980 3206 5000 3210
rect 4800 3150 4820 3154
rect 4880 3150 4920 3154
rect 4980 3150 5000 3154
rect 4800 3140 5000 3150
rect 6000 3210 6200 3220
rect 6000 3206 6020 3210
rect 6080 3206 6120 3210
rect 6180 3206 6200 3210
rect 6000 3150 6020 3154
rect 6080 3150 6120 3154
rect 6180 3150 6200 3154
rect 6000 3140 6200 3150
rect 7200 3210 7400 3220
rect 7200 3206 7220 3210
rect 7280 3206 7320 3210
rect 7380 3206 7400 3210
rect 7200 3150 7220 3154
rect 7280 3150 7320 3154
rect 7380 3150 7400 3154
rect 7200 3140 7400 3150
rect 8400 3210 8600 3220
rect 8400 3206 8420 3210
rect 8480 3206 8520 3210
rect 8580 3206 8600 3210
rect 8400 3150 8420 3154
rect 8480 3150 8520 3154
rect 8580 3150 8600 3154
rect 8400 3140 8600 3150
rect 9600 3210 9800 3220
rect 9600 3206 9620 3210
rect 9680 3206 9720 3210
rect 9780 3206 9800 3210
rect 9600 3150 9620 3154
rect 9680 3150 9720 3154
rect 9780 3150 9800 3154
rect 9600 3140 9800 3150
rect 10800 3210 11000 3220
rect 10800 3206 10820 3210
rect 10880 3206 10920 3210
rect 10980 3206 11000 3210
rect 10800 3150 10820 3154
rect 10880 3150 10920 3154
rect 10980 3150 11000 3154
rect 10800 3140 11000 3150
rect 12000 3210 12200 3220
rect 12000 3206 12020 3210
rect 12080 3206 12120 3210
rect 12180 3206 12200 3210
rect 12000 3150 12020 3154
rect 12080 3150 12120 3154
rect 12180 3150 12200 3154
rect 12000 3140 12200 3150
rect 13200 3210 13400 3220
rect 13200 3206 13220 3210
rect 13280 3206 13320 3210
rect 13380 3206 13400 3210
rect 13200 3150 13220 3154
rect 13280 3150 13320 3154
rect 13380 3150 13400 3154
rect 13200 3140 13400 3150
rect 14400 3210 14600 3220
rect 14400 3206 14420 3210
rect 14480 3206 14520 3210
rect 14580 3206 14600 3210
rect 14400 3150 14420 3154
rect 14480 3150 14520 3154
rect 14580 3150 14600 3154
rect 14400 3140 14600 3150
rect 15600 3210 15800 3220
rect 15600 3206 15620 3210
rect 15680 3206 15720 3210
rect 15780 3206 15800 3210
rect 15600 3150 15620 3154
rect 15680 3150 15720 3154
rect 15780 3150 15800 3154
rect 15600 3140 15800 3150
rect 16800 3210 17000 3220
rect 16800 3206 16820 3210
rect 16880 3206 16920 3210
rect 16980 3206 17000 3210
rect 16800 3150 16820 3154
rect 16880 3150 16920 3154
rect 16980 3150 17000 3154
rect 16800 3140 17000 3150
rect 18000 3210 18200 3220
rect 18000 3206 18020 3210
rect 18080 3206 18120 3210
rect 18180 3206 18200 3210
rect 18000 3150 18020 3154
rect 18080 3150 18120 3154
rect 18180 3150 18200 3154
rect 18000 3140 18200 3150
rect 19200 3210 19400 3220
rect 19200 3206 19220 3210
rect 19280 3206 19320 3210
rect 19380 3206 19400 3210
rect 19200 3150 19220 3154
rect 19280 3150 19320 3154
rect 19380 3150 19400 3154
rect 19200 3140 19400 3150
rect 0 2814 200 2824
rect 0 2810 20 2814
rect 80 2810 120 2814
rect 180 2810 200 2814
rect 0 2754 20 2758
rect 80 2754 120 2758
rect 180 2754 200 2758
rect 0 2744 200 2754
rect 1200 2814 1400 2824
rect 1200 2810 1220 2814
rect 1280 2810 1320 2814
rect 1380 2810 1400 2814
rect 1200 2754 1220 2758
rect 1280 2754 1320 2758
rect 1380 2754 1400 2758
rect 1200 2744 1400 2754
rect 2400 2814 2600 2824
rect 2400 2810 2420 2814
rect 2480 2810 2520 2814
rect 2580 2810 2600 2814
rect 2400 2754 2420 2758
rect 2480 2754 2520 2758
rect 2580 2754 2600 2758
rect 2400 2744 2600 2754
rect 3600 2814 3800 2824
rect 3600 2810 3620 2814
rect 3680 2810 3720 2814
rect 3780 2810 3800 2814
rect 3600 2754 3620 2758
rect 3680 2754 3720 2758
rect 3780 2754 3800 2758
rect 3600 2744 3800 2754
rect 4800 2814 5000 2824
rect 4800 2810 4820 2814
rect 4880 2810 4920 2814
rect 4980 2810 5000 2814
rect 4800 2754 4820 2758
rect 4880 2754 4920 2758
rect 4980 2754 5000 2758
rect 4800 2744 5000 2754
rect 6000 2814 6200 2824
rect 6000 2810 6020 2814
rect 6080 2810 6120 2814
rect 6180 2810 6200 2814
rect 6000 2754 6020 2758
rect 6080 2754 6120 2758
rect 6180 2754 6200 2758
rect 6000 2744 6200 2754
rect 7200 2814 7400 2824
rect 7200 2810 7220 2814
rect 7280 2810 7320 2814
rect 7380 2810 7400 2814
rect 7200 2754 7220 2758
rect 7280 2754 7320 2758
rect 7380 2754 7400 2758
rect 7200 2744 7400 2754
rect 8400 2814 8600 2824
rect 8400 2810 8420 2814
rect 8480 2810 8520 2814
rect 8580 2810 8600 2814
rect 8400 2754 8420 2758
rect 8480 2754 8520 2758
rect 8580 2754 8600 2758
rect 8400 2744 8600 2754
rect 9600 2814 9800 2824
rect 9600 2810 9620 2814
rect 9680 2810 9720 2814
rect 9780 2810 9800 2814
rect 9600 2754 9620 2758
rect 9680 2754 9720 2758
rect 9780 2754 9800 2758
rect 9600 2744 9800 2754
rect 10800 2814 11000 2824
rect 10800 2810 10820 2814
rect 10880 2810 10920 2814
rect 10980 2810 11000 2814
rect 10800 2754 10820 2758
rect 10880 2754 10920 2758
rect 10980 2754 11000 2758
rect 10800 2744 11000 2754
rect 12000 2814 12200 2824
rect 12000 2810 12020 2814
rect 12080 2810 12120 2814
rect 12180 2810 12200 2814
rect 12000 2754 12020 2758
rect 12080 2754 12120 2758
rect 12180 2754 12200 2758
rect 12000 2744 12200 2754
rect 13200 2814 13400 2824
rect 13200 2810 13220 2814
rect 13280 2810 13320 2814
rect 13380 2810 13400 2814
rect 13200 2754 13220 2758
rect 13280 2754 13320 2758
rect 13380 2754 13400 2758
rect 13200 2744 13400 2754
rect 14400 2814 14600 2824
rect 14400 2810 14420 2814
rect 14480 2810 14520 2814
rect 14580 2810 14600 2814
rect 14400 2754 14420 2758
rect 14480 2754 14520 2758
rect 14580 2754 14600 2758
rect 14400 2744 14600 2754
rect 15600 2814 15800 2824
rect 15600 2810 15620 2814
rect 15680 2810 15720 2814
rect 15780 2810 15800 2814
rect 15600 2754 15620 2758
rect 15680 2754 15720 2758
rect 15780 2754 15800 2758
rect 15600 2744 15800 2754
rect 16800 2814 17000 2824
rect 16800 2810 16820 2814
rect 16880 2810 16920 2814
rect 16980 2810 17000 2814
rect 16800 2754 16820 2758
rect 16880 2754 16920 2758
rect 16980 2754 17000 2758
rect 16800 2744 17000 2754
rect 18000 2814 18200 2824
rect 18000 2810 18020 2814
rect 18080 2810 18120 2814
rect 18180 2810 18200 2814
rect 18000 2754 18020 2758
rect 18080 2754 18120 2758
rect 18180 2754 18200 2758
rect 18000 2744 18200 2754
rect 19200 2814 19400 2824
rect 19200 2810 19220 2814
rect 19280 2810 19320 2814
rect 19380 2810 19400 2814
rect 19200 2754 19220 2758
rect 19280 2754 19320 2758
rect 19380 2754 19400 2758
rect 19200 2744 19400 2754
rect 20400 2814 20600 2824
rect 20400 2810 20420 2814
rect 20480 2810 20520 2814
rect 20580 2810 20600 2814
rect 20400 2754 20420 2758
rect 20480 2754 20520 2758
rect 20580 2754 20600 2758
rect 20400 2744 20600 2754
rect 21156 2814 21356 2824
rect 21156 2810 21176 2814
rect 21236 2810 21276 2814
rect 21336 2810 21356 2814
rect 21156 2754 21176 2758
rect 21236 2754 21276 2758
rect 21336 2754 21356 2758
rect 21156 2744 21356 2754
<< via2 >>
rect 20408 3888 20488 3894
rect 20408 3820 20414 3888
rect 20414 3820 20482 3888
rect 20482 3820 20488 3888
rect 20408 3814 20488 3820
rect 20512 3888 20592 3894
rect 20512 3820 20518 3888
rect 20518 3820 20586 3888
rect 20586 3820 20592 3888
rect 20512 3814 20592 3820
rect 20408 3784 20488 3790
rect 20408 3716 20414 3784
rect 20414 3716 20482 3784
rect 20482 3716 20488 3784
rect 20408 3710 20488 3716
rect 20512 3784 20592 3790
rect 20512 3716 20518 3784
rect 20518 3716 20586 3784
rect 20586 3716 20592 3784
rect 20512 3710 20592 3716
rect 2420 3206 2480 3210
rect 2520 3206 2580 3210
rect 2420 3154 2452 3206
rect 2452 3154 2474 3206
rect 2474 3154 2480 3206
rect 2520 3154 2526 3206
rect 2526 3154 2548 3206
rect 2548 3154 2580 3206
rect 2420 3150 2480 3154
rect 2520 3150 2580 3154
rect 3620 3206 3680 3210
rect 3720 3206 3780 3210
rect 3620 3154 3652 3206
rect 3652 3154 3674 3206
rect 3674 3154 3680 3206
rect 3720 3154 3726 3206
rect 3726 3154 3748 3206
rect 3748 3154 3780 3206
rect 3620 3150 3680 3154
rect 3720 3150 3780 3154
rect 4820 3206 4880 3210
rect 4920 3206 4980 3210
rect 4820 3154 4852 3206
rect 4852 3154 4874 3206
rect 4874 3154 4880 3206
rect 4920 3154 4926 3206
rect 4926 3154 4948 3206
rect 4948 3154 4980 3206
rect 4820 3150 4880 3154
rect 4920 3150 4980 3154
rect 6020 3206 6080 3210
rect 6120 3206 6180 3210
rect 6020 3154 6052 3206
rect 6052 3154 6074 3206
rect 6074 3154 6080 3206
rect 6120 3154 6126 3206
rect 6126 3154 6148 3206
rect 6148 3154 6180 3206
rect 6020 3150 6080 3154
rect 6120 3150 6180 3154
rect 7220 3206 7280 3210
rect 7320 3206 7380 3210
rect 7220 3154 7252 3206
rect 7252 3154 7274 3206
rect 7274 3154 7280 3206
rect 7320 3154 7326 3206
rect 7326 3154 7348 3206
rect 7348 3154 7380 3206
rect 7220 3150 7280 3154
rect 7320 3150 7380 3154
rect 8420 3206 8480 3210
rect 8520 3206 8580 3210
rect 8420 3154 8452 3206
rect 8452 3154 8474 3206
rect 8474 3154 8480 3206
rect 8520 3154 8526 3206
rect 8526 3154 8548 3206
rect 8548 3154 8580 3206
rect 8420 3150 8480 3154
rect 8520 3150 8580 3154
rect 9620 3206 9680 3210
rect 9720 3206 9780 3210
rect 9620 3154 9652 3206
rect 9652 3154 9674 3206
rect 9674 3154 9680 3206
rect 9720 3154 9726 3206
rect 9726 3154 9748 3206
rect 9748 3154 9780 3206
rect 9620 3150 9680 3154
rect 9720 3150 9780 3154
rect 10820 3206 10880 3210
rect 10920 3206 10980 3210
rect 10820 3154 10852 3206
rect 10852 3154 10874 3206
rect 10874 3154 10880 3206
rect 10920 3154 10926 3206
rect 10926 3154 10948 3206
rect 10948 3154 10980 3206
rect 10820 3150 10880 3154
rect 10920 3150 10980 3154
rect 12020 3206 12080 3210
rect 12120 3206 12180 3210
rect 12020 3154 12052 3206
rect 12052 3154 12074 3206
rect 12074 3154 12080 3206
rect 12120 3154 12126 3206
rect 12126 3154 12148 3206
rect 12148 3154 12180 3206
rect 12020 3150 12080 3154
rect 12120 3150 12180 3154
rect 13220 3206 13280 3210
rect 13320 3206 13380 3210
rect 13220 3154 13252 3206
rect 13252 3154 13274 3206
rect 13274 3154 13280 3206
rect 13320 3154 13326 3206
rect 13326 3154 13348 3206
rect 13348 3154 13380 3206
rect 13220 3150 13280 3154
rect 13320 3150 13380 3154
rect 14420 3206 14480 3210
rect 14520 3206 14580 3210
rect 14420 3154 14452 3206
rect 14452 3154 14474 3206
rect 14474 3154 14480 3206
rect 14520 3154 14526 3206
rect 14526 3154 14548 3206
rect 14548 3154 14580 3206
rect 14420 3150 14480 3154
rect 14520 3150 14580 3154
rect 15620 3206 15680 3210
rect 15720 3206 15780 3210
rect 15620 3154 15652 3206
rect 15652 3154 15674 3206
rect 15674 3154 15680 3206
rect 15720 3154 15726 3206
rect 15726 3154 15748 3206
rect 15748 3154 15780 3206
rect 15620 3150 15680 3154
rect 15720 3150 15780 3154
rect 16820 3206 16880 3210
rect 16920 3206 16980 3210
rect 16820 3154 16852 3206
rect 16852 3154 16874 3206
rect 16874 3154 16880 3206
rect 16920 3154 16926 3206
rect 16926 3154 16948 3206
rect 16948 3154 16980 3206
rect 16820 3150 16880 3154
rect 16920 3150 16980 3154
rect 18020 3206 18080 3210
rect 18120 3206 18180 3210
rect 18020 3154 18052 3206
rect 18052 3154 18074 3206
rect 18074 3154 18080 3206
rect 18120 3154 18126 3206
rect 18126 3154 18148 3206
rect 18148 3154 18180 3206
rect 18020 3150 18080 3154
rect 18120 3150 18180 3154
rect 19220 3206 19280 3210
rect 19320 3206 19380 3210
rect 19220 3154 19252 3206
rect 19252 3154 19274 3206
rect 19274 3154 19280 3206
rect 19320 3154 19326 3206
rect 19326 3154 19348 3206
rect 19348 3154 19380 3206
rect 19220 3150 19280 3154
rect 19320 3150 19380 3154
rect 20 2810 80 2814
rect 120 2810 180 2814
rect 20 2758 52 2810
rect 52 2758 74 2810
rect 74 2758 80 2810
rect 120 2758 126 2810
rect 126 2758 148 2810
rect 148 2758 180 2810
rect 20 2754 80 2758
rect 120 2754 180 2758
rect 1220 2810 1280 2814
rect 1320 2810 1380 2814
rect 1220 2758 1252 2810
rect 1252 2758 1274 2810
rect 1274 2758 1280 2810
rect 1320 2758 1326 2810
rect 1326 2758 1348 2810
rect 1348 2758 1380 2810
rect 1220 2754 1280 2758
rect 1320 2754 1380 2758
rect 2420 2810 2480 2814
rect 2520 2810 2580 2814
rect 2420 2758 2452 2810
rect 2452 2758 2474 2810
rect 2474 2758 2480 2810
rect 2520 2758 2526 2810
rect 2526 2758 2548 2810
rect 2548 2758 2580 2810
rect 2420 2754 2480 2758
rect 2520 2754 2580 2758
rect 3620 2810 3680 2814
rect 3720 2810 3780 2814
rect 3620 2758 3652 2810
rect 3652 2758 3674 2810
rect 3674 2758 3680 2810
rect 3720 2758 3726 2810
rect 3726 2758 3748 2810
rect 3748 2758 3780 2810
rect 3620 2754 3680 2758
rect 3720 2754 3780 2758
rect 4820 2810 4880 2814
rect 4920 2810 4980 2814
rect 4820 2758 4852 2810
rect 4852 2758 4874 2810
rect 4874 2758 4880 2810
rect 4920 2758 4926 2810
rect 4926 2758 4948 2810
rect 4948 2758 4980 2810
rect 4820 2754 4880 2758
rect 4920 2754 4980 2758
rect 6020 2810 6080 2814
rect 6120 2810 6180 2814
rect 6020 2758 6052 2810
rect 6052 2758 6074 2810
rect 6074 2758 6080 2810
rect 6120 2758 6126 2810
rect 6126 2758 6148 2810
rect 6148 2758 6180 2810
rect 6020 2754 6080 2758
rect 6120 2754 6180 2758
rect 7220 2810 7280 2814
rect 7320 2810 7380 2814
rect 7220 2758 7252 2810
rect 7252 2758 7274 2810
rect 7274 2758 7280 2810
rect 7320 2758 7326 2810
rect 7326 2758 7348 2810
rect 7348 2758 7380 2810
rect 7220 2754 7280 2758
rect 7320 2754 7380 2758
rect 8420 2810 8480 2814
rect 8520 2810 8580 2814
rect 8420 2758 8452 2810
rect 8452 2758 8474 2810
rect 8474 2758 8480 2810
rect 8520 2758 8526 2810
rect 8526 2758 8548 2810
rect 8548 2758 8580 2810
rect 8420 2754 8480 2758
rect 8520 2754 8580 2758
rect 9620 2810 9680 2814
rect 9720 2810 9780 2814
rect 9620 2758 9652 2810
rect 9652 2758 9674 2810
rect 9674 2758 9680 2810
rect 9720 2758 9726 2810
rect 9726 2758 9748 2810
rect 9748 2758 9780 2810
rect 9620 2754 9680 2758
rect 9720 2754 9780 2758
rect 10820 2810 10880 2814
rect 10920 2810 10980 2814
rect 10820 2758 10852 2810
rect 10852 2758 10874 2810
rect 10874 2758 10880 2810
rect 10920 2758 10926 2810
rect 10926 2758 10948 2810
rect 10948 2758 10980 2810
rect 10820 2754 10880 2758
rect 10920 2754 10980 2758
rect 12020 2810 12080 2814
rect 12120 2810 12180 2814
rect 12020 2758 12052 2810
rect 12052 2758 12074 2810
rect 12074 2758 12080 2810
rect 12120 2758 12126 2810
rect 12126 2758 12148 2810
rect 12148 2758 12180 2810
rect 12020 2754 12080 2758
rect 12120 2754 12180 2758
rect 13220 2810 13280 2814
rect 13320 2810 13380 2814
rect 13220 2758 13252 2810
rect 13252 2758 13274 2810
rect 13274 2758 13280 2810
rect 13320 2758 13326 2810
rect 13326 2758 13348 2810
rect 13348 2758 13380 2810
rect 13220 2754 13280 2758
rect 13320 2754 13380 2758
rect 14420 2810 14480 2814
rect 14520 2810 14580 2814
rect 14420 2758 14452 2810
rect 14452 2758 14474 2810
rect 14474 2758 14480 2810
rect 14520 2758 14526 2810
rect 14526 2758 14548 2810
rect 14548 2758 14580 2810
rect 14420 2754 14480 2758
rect 14520 2754 14580 2758
rect 15620 2810 15680 2814
rect 15720 2810 15780 2814
rect 15620 2758 15652 2810
rect 15652 2758 15674 2810
rect 15674 2758 15680 2810
rect 15720 2758 15726 2810
rect 15726 2758 15748 2810
rect 15748 2758 15780 2810
rect 15620 2754 15680 2758
rect 15720 2754 15780 2758
rect 16820 2810 16880 2814
rect 16920 2810 16980 2814
rect 16820 2758 16852 2810
rect 16852 2758 16874 2810
rect 16874 2758 16880 2810
rect 16920 2758 16926 2810
rect 16926 2758 16948 2810
rect 16948 2758 16980 2810
rect 16820 2754 16880 2758
rect 16920 2754 16980 2758
rect 18020 2810 18080 2814
rect 18120 2810 18180 2814
rect 18020 2758 18052 2810
rect 18052 2758 18074 2810
rect 18074 2758 18080 2810
rect 18120 2758 18126 2810
rect 18126 2758 18148 2810
rect 18148 2758 18180 2810
rect 18020 2754 18080 2758
rect 18120 2754 18180 2758
rect 19220 2810 19280 2814
rect 19320 2810 19380 2814
rect 19220 2758 19252 2810
rect 19252 2758 19274 2810
rect 19274 2758 19280 2810
rect 19320 2758 19326 2810
rect 19326 2758 19348 2810
rect 19348 2758 19380 2810
rect 19220 2754 19280 2758
rect 19320 2754 19380 2758
rect 20420 2810 20480 2814
rect 20520 2810 20580 2814
rect 20420 2758 20452 2810
rect 20452 2758 20474 2810
rect 20474 2758 20480 2810
rect 20520 2758 20526 2810
rect 20526 2758 20548 2810
rect 20548 2758 20580 2810
rect 20420 2754 20480 2758
rect 20520 2754 20580 2758
rect 21176 2810 21236 2814
rect 21276 2810 21336 2814
rect 21176 2758 21208 2810
rect 21208 2758 21230 2810
rect 21230 2758 21236 2810
rect 21276 2758 21282 2810
rect 21282 2758 21304 2810
rect 21304 2758 21336 2810
rect 21176 2754 21236 2758
rect 21276 2754 21336 2758
<< metal3 >>
rect 20400 3894 20600 3903
rect 20400 3814 20408 3894
rect 20488 3814 20512 3894
rect 20592 3814 20600 3894
rect 20400 3790 20600 3814
rect 20400 3710 20408 3790
rect 20488 3710 20512 3790
rect 20592 3710 20600 3790
rect 2400 3210 2600 3230
rect 2400 3150 2420 3210
rect 2480 3150 2520 3210
rect 2580 3150 2600 3210
rect 2400 3134 2600 3150
rect 3600 3210 3800 3230
rect 3600 3150 3620 3210
rect 3680 3150 3720 3210
rect 3780 3150 3800 3210
rect 3600 3134 3800 3150
rect 4800 3210 5000 3230
rect 4800 3150 4820 3210
rect 4880 3150 4920 3210
rect 4980 3150 5000 3210
rect 4800 3134 5000 3150
rect 6000 3210 6200 3230
rect 6000 3150 6020 3210
rect 6080 3150 6120 3210
rect 6180 3150 6200 3210
rect 6000 3134 6200 3150
rect 7200 3210 7400 3230
rect 7200 3150 7220 3210
rect 7280 3150 7320 3210
rect 7380 3150 7400 3210
rect 7200 3134 7400 3150
rect 8400 3210 8600 3230
rect 8400 3150 8420 3210
rect 8480 3150 8520 3210
rect 8580 3150 8600 3210
rect 8400 3134 8600 3150
rect 9600 3210 9800 3230
rect 9600 3150 9620 3210
rect 9680 3150 9720 3210
rect 9780 3150 9800 3210
rect 9600 3134 9800 3150
rect 10800 3210 11000 3230
rect 10800 3150 10820 3210
rect 10880 3150 10920 3210
rect 10980 3150 11000 3210
rect 10800 3134 11000 3150
rect 12000 3210 12200 3230
rect 12000 3150 12020 3210
rect 12080 3150 12120 3210
rect 12180 3150 12200 3210
rect 12000 3134 12200 3150
rect 13200 3210 13400 3230
rect 13200 3150 13220 3210
rect 13280 3150 13320 3210
rect 13380 3150 13400 3210
rect 13200 3134 13400 3150
rect 14400 3210 14600 3230
rect 14400 3150 14420 3210
rect 14480 3150 14520 3210
rect 14580 3150 14600 3210
rect 14400 3134 14600 3150
rect 15600 3210 15800 3230
rect 15600 3150 15620 3210
rect 15680 3150 15720 3210
rect 15780 3150 15800 3210
rect 15600 3134 15800 3150
rect 16800 3210 17000 3230
rect 16800 3150 16820 3210
rect 16880 3150 16920 3210
rect 16980 3150 17000 3210
rect 16800 3134 17000 3150
rect 18000 3210 18200 3230
rect 18000 3150 18020 3210
rect 18080 3150 18120 3210
rect 18180 3150 18200 3210
rect 18000 3134 18200 3150
rect 19200 3210 19400 3230
rect 19200 3150 19220 3210
rect 19280 3150 19320 3210
rect 19380 3150 19400 3210
rect 19200 3134 19400 3150
rect 20400 3134 20600 3710
rect 0 2834 21356 3134
rect 0 2814 200 2834
rect 0 2754 20 2814
rect 80 2754 120 2814
rect 180 2754 200 2814
rect 0 2738 200 2754
rect 1200 2814 1400 2834
rect 1200 2754 1220 2814
rect 1280 2754 1320 2814
rect 1380 2754 1400 2814
rect 1200 2738 1400 2754
rect 2400 2814 2600 2834
rect 2400 2754 2420 2814
rect 2480 2754 2520 2814
rect 2580 2754 2600 2814
rect 2400 2738 2600 2754
rect 3600 2814 3800 2834
rect 3600 2754 3620 2814
rect 3680 2754 3720 2814
rect 3780 2754 3800 2814
rect 3600 2738 3800 2754
rect 4800 2814 5000 2834
rect 4800 2754 4820 2814
rect 4880 2754 4920 2814
rect 4980 2754 5000 2814
rect 4800 2738 5000 2754
rect 6000 2814 6200 2834
rect 6000 2754 6020 2814
rect 6080 2754 6120 2814
rect 6180 2754 6200 2814
rect 6000 2738 6200 2754
rect 7200 2814 7400 2834
rect 7200 2754 7220 2814
rect 7280 2754 7320 2814
rect 7380 2754 7400 2814
rect 7200 2738 7400 2754
rect 8400 2814 8600 2834
rect 8400 2754 8420 2814
rect 8480 2754 8520 2814
rect 8580 2754 8600 2814
rect 8400 2738 8600 2754
rect 9600 2814 9800 2834
rect 9600 2754 9620 2814
rect 9680 2754 9720 2814
rect 9780 2754 9800 2814
rect 9600 2738 9800 2754
rect 10800 2814 11000 2834
rect 10800 2754 10820 2814
rect 10880 2754 10920 2814
rect 10980 2754 11000 2814
rect 10800 2738 11000 2754
rect 12000 2814 12200 2834
rect 12000 2754 12020 2814
rect 12080 2754 12120 2814
rect 12180 2754 12200 2814
rect 12000 2738 12200 2754
rect 13200 2814 13400 2834
rect 13200 2754 13220 2814
rect 13280 2754 13320 2814
rect 13380 2754 13400 2814
rect 13200 2738 13400 2754
rect 14400 2814 14600 2834
rect 14400 2754 14420 2814
rect 14480 2754 14520 2814
rect 14580 2754 14600 2814
rect 14400 2738 14600 2754
rect 15600 2814 15800 2834
rect 15600 2754 15620 2814
rect 15680 2754 15720 2814
rect 15780 2754 15800 2814
rect 15600 2738 15800 2754
rect 16800 2814 17000 2834
rect 16800 2754 16820 2814
rect 16880 2754 16920 2814
rect 16980 2754 17000 2814
rect 16800 2738 17000 2754
rect 18000 2814 18200 2834
rect 18000 2754 18020 2814
rect 18080 2754 18120 2814
rect 18180 2754 18200 2814
rect 18000 2738 18200 2754
rect 19200 2814 19400 2834
rect 19200 2754 19220 2814
rect 19280 2754 19320 2814
rect 19380 2754 19400 2814
rect 19200 2738 19400 2754
rect 20400 2814 20600 2834
rect 20400 2754 20420 2814
rect 20480 2754 20520 2814
rect 20580 2754 20600 2814
rect 20400 2738 20600 2754
rect 21156 2814 21356 2834
rect 21156 2754 21176 2814
rect 21236 2754 21276 2814
rect 21336 2754 21356 2814
rect 21156 2738 21356 2754
use inv  inv_5
timestamp 1623637110
transform -1 0 3246 0 -1 4834
box -400 1960 3246 4834
use inv  inv_4
timestamp 1623637110
transform -1 0 6788 0 -1 4834
box -400 1960 3246 4834
use inv  inv_3
timestamp 1623637110
transform -1 0 10330 0 -1 4834
box -400 1960 3246 4834
use inv  inv_2
timestamp 1623637110
transform -1 0 13872 0 -1 4834
box -400 1960 3246 4834
use inv  inv_1
timestamp 1623637110
transform -1 0 17414 0 -1 4834
box -400 1960 3246 4834
use inv  inv_0
timestamp 1623637110
transform -1 0 20956 0 -1 4834
box -400 1960 3246 4834
use inv  inv_6
timestamp 1623637110
transform 1 0 2096 0 1 1134
box -400 1960 3246 4834
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621367673
transform 1 0 637 0 1 4560
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621367673
transform 1 0 -162 0 1 4560
box -38 -48 498 592
use inv  inv_7
timestamp 1623637110
transform 1 0 5638 0 1 1134
box -400 1960 3246 4834
use inv  inv_8
timestamp 1623637110
transform 1 0 9180 0 1 1134
box -400 1960 3246 4834
use inv  inv_9
timestamp 1623637110
transform 1 0 12722 0 1 1134
box -400 1960 3246 4834
use inv  inv_10
timestamp 1623637110
transform 1 0 16264 0 1 1134
box -400 1960 3246 4834
use res_poly  res_poly_0
timestamp 1623640090
transform 1 0 20200 0 1 3900
box -100 -100 500 1100
use res_poly  res_poly_1
timestamp 1623640090
transform 0 1 20600 -1 0 3900
box -100 -100 500 1100
<< labels >>
flabel metal1 17728 1106 17800 1178 1 FreeSans 200 0 0 0 p[0]  
flabel metal1 14182 1106 14254 1178 1 FreeSans 200 0 0 0 p[1]        
flabel metal1 10650 1106 10722 1178 1 FreeSans 200 0 0 0 p[2]        
flabel metal1 7106 1106 7178 1178 1 FreeSans 200 0 0 0 p[3]
flabel metal1 3556 1106 3628 1178 1 FreeSans 200 0 0 0 p[4]
flabel metal1 -72 1106 0 1178 1 FreeSans 200 0 0 0 p[5]
flabel metal1 5254 4790 5326 4862 1 FreeSans 200 0 0 0 p[6]
flabel metal1 8796 4790 8868 4862 1 FreeSans 200 0 0 0 p[7]
flabel metal1 12334 4790 12406 4862 1 FreeSans 200 0 0 0 p[8]
flabel metal1 15878 4790 15950 4862 1 FreeSans 200 0 0 0 p[9]
flabel metal1 19510 4790 19582 4862 1 FreeSans 200 0 0 0 p[10]
flabel metal1 17728 1650 17800 1722 1 FreeSans 200 0 0 0 pn[0]
flabel metal1 14182 1650 14254 1722 1 FreeSans 200 0 0 0 pn[1]
flabel metal1 10634 1650 10706 1722 1 FreeSans 200 0 0 0 pn[2]
flabel metal1 7104 1650 7176 1722 1 FreeSans 200 0 0 0 pn[3]
flabel metal1 3554 1650 3626 1722 1 FreeSans 200 0 0 0 pn[4]
flabel metal1 -72 1650 0 1722 1 FreeSans 200 0 0 0 pn[5]
flabel metal1 5254 4246 5326 4318 1 FreeSans 200 0 0 0 pn[6]
flabel metal1 8798 4246 8870 4318 1 FreeSans 200 0 0 0 pn[7]
flabel metal1 12334 4246 12406 4318 1 FreeSans 200 0 0 0 pn[8]
flabel metal1 15878 4246 15950 4318 1 FreeSans 200 0 0 0 pn[9]
flabel metal1 19510 4246 19582 4318 1 FreeSans 200 0 0 0 pn[10]
flabel metal2 21600 3800 21700 3900 1 FreeSans 200 0 0 0 input_analog
flabel metal3 20400 3498 20502 3600 1 FreeSans 200 0 0 0 v_ctr
flabel metal1 -200 4512 -104 4608 1 FreeSans 200 0 0 0 vssd2
flabel metal1 -200 5056 -104 5152 1 FreeSans 200 0 0 0 vccd2
flabel metal1 1680 5854 1776 5950 1 FreeSans 200 0 0 0 vccd2
flabel metal1 20524 4804 20596 4876 1 FreeSans 200 0 0 0 vssd2
<< end >>
