magic
tech sky130A
magscale 1 2
timestamp 1637941551
<< poly >>
rect 0 955 400 976
rect 0 921 22 955
rect 56 921 102 955
rect 136 921 182 955
rect 216 921 262 955
rect 296 921 342 955
rect 376 921 400 955
rect 0 903 400 921
rect 0 52 400 73
rect 0 18 22 52
rect 56 18 102 52
rect 136 18 182 52
rect 216 18 262 52
rect 296 18 342 52
rect 376 18 400 52
rect 0 -6 400 18
<< polycont >>
rect 22 921 56 955
rect 102 921 136 955
rect 182 921 216 955
rect 262 921 296 955
rect 342 921 376 955
rect 22 18 56 52
rect 102 18 136 52
rect 182 18 216 52
rect 262 18 296 52
rect 342 18 376 52
<< npolyres >>
rect 0 73 400 903
<< locali >>
rect 0 955 400 976
rect 0 921 22 955
rect 56 921 102 955
rect 136 921 182 955
rect 216 921 262 955
rect 296 921 342 955
rect 376 921 400 955
rect 0 903 400 921
rect 0 52 400 73
rect 0 18 22 52
rect 56 18 102 52
rect 136 18 182 52
rect 216 18 262 52
rect 296 18 342 52
rect 376 18 400 52
rect 0 0 400 18
<< end >>
