magic
tech sky130A
timestamp 1637172953
<< pwell >>
rect 0 0 400 610
<< nmos >>
rect 105 100 295 500
<< ndiff >>
rect 75 489 105 500
rect 75 471 81 489
rect 99 471 105 489
rect 75 453 105 471
rect 75 435 81 453
rect 99 435 105 453
rect 75 417 105 435
rect 75 399 81 417
rect 99 399 105 417
rect 75 381 105 399
rect 75 363 81 381
rect 99 363 105 381
rect 75 345 105 363
rect 75 327 81 345
rect 99 327 105 345
rect 75 309 105 327
rect 75 291 81 309
rect 99 291 105 309
rect 75 273 105 291
rect 75 255 81 273
rect 99 255 105 273
rect 75 237 105 255
rect 75 219 81 237
rect 99 219 105 237
rect 75 201 105 219
rect 75 183 81 201
rect 99 183 105 201
rect 75 165 105 183
rect 75 147 81 165
rect 99 147 105 165
rect 75 129 105 147
rect 75 111 81 129
rect 99 111 105 129
rect 75 100 105 111
rect 295 489 325 500
rect 295 471 301 489
rect 319 471 325 489
rect 295 453 325 471
rect 295 435 301 453
rect 319 435 325 453
rect 295 417 325 435
rect 295 399 301 417
rect 319 399 325 417
rect 295 381 325 399
rect 295 363 301 381
rect 319 363 325 381
rect 295 345 325 363
rect 295 327 301 345
rect 319 327 325 345
rect 295 309 325 327
rect 295 291 301 309
rect 319 291 325 309
rect 295 273 325 291
rect 295 255 301 273
rect 319 255 325 273
rect 295 237 325 255
rect 295 219 301 237
rect 319 219 325 237
rect 295 201 325 219
rect 295 183 301 201
rect 319 183 325 201
rect 295 165 325 183
rect 295 147 301 165
rect 319 147 325 165
rect 295 129 325 147
rect 295 111 301 129
rect 319 111 325 129
rect 295 100 325 111
<< ndiffc >>
rect 81 471 99 489
rect 81 435 99 453
rect 81 399 99 417
rect 81 363 99 381
rect 81 327 99 345
rect 81 291 99 309
rect 81 255 99 273
rect 81 219 99 237
rect 81 183 99 201
rect 81 147 99 165
rect 81 111 99 129
rect 301 471 319 489
rect 301 435 319 453
rect 301 399 319 417
rect 301 363 319 381
rect 301 327 319 345
rect 301 291 319 309
rect 301 255 319 273
rect 301 219 319 237
rect 301 183 319 201
rect 301 147 319 165
rect 301 111 319 129
<< poly >>
rect 105 500 295 544
rect 105 87 295 100
<< locali >>
rect 75 489 105 502
rect 75 471 81 489
rect 99 471 105 489
rect 75 453 105 471
rect 75 435 81 453
rect 99 435 105 453
rect 75 417 105 435
rect 75 399 81 417
rect 99 399 105 417
rect 75 381 105 399
rect 75 363 81 381
rect 99 363 105 381
rect 75 345 105 363
rect 75 327 81 345
rect 99 327 105 345
rect 75 309 105 327
rect 75 291 81 309
rect 99 291 105 309
rect 75 273 105 291
rect 75 255 81 273
rect 99 255 105 273
rect 75 237 105 255
rect 75 219 81 237
rect 99 219 105 237
rect 75 201 105 219
rect 75 183 81 201
rect 99 183 105 201
rect 75 165 105 183
rect 75 147 81 165
rect 99 147 105 165
rect 75 129 105 147
rect 75 111 81 129
rect 99 111 105 129
rect 75 98 105 111
rect 295 489 325 502
rect 295 471 301 489
rect 319 471 325 489
rect 295 453 325 471
rect 295 435 301 453
rect 319 435 325 453
rect 295 417 325 435
rect 295 399 301 417
rect 319 399 325 417
rect 295 381 325 399
rect 295 363 301 381
rect 319 363 325 381
rect 295 345 325 363
rect 295 327 301 345
rect 319 327 325 345
rect 295 309 325 327
rect 295 291 301 309
rect 319 291 325 309
rect 295 273 325 291
rect 295 255 301 273
rect 319 255 325 273
rect 295 237 325 255
rect 295 219 301 237
rect 319 219 325 237
rect 295 201 325 219
rect 295 183 301 201
rect 319 183 325 201
rect 295 165 325 183
rect 295 147 301 165
rect 319 147 325 165
rect 295 129 325 147
rect 295 111 301 129
rect 319 111 325 129
rect 295 98 325 111
<< end >>
