magic
tech sky130A
timestamp 1637401559
<< metal1 >>
rect 300 2553 652 2603
rect 8973 2553 9450 2603
rect 300 2000 350 2553
rect -300 1950 350 2000
rect 450 2253 602 2303
rect 9153 2253 9300 2303
rect -300 885 -250 1950
rect 450 1850 500 2253
rect -150 1800 500 1850
rect 603 1859 703 1866
rect 603 1829 610 1859
rect 640 1829 666 1859
rect 696 1829 703 1859
rect 603 1822 703 1829
rect 1051 1859 1263 1866
rect 1051 1829 1058 1859
rect 1088 1829 1114 1859
rect 1144 1829 1170 1859
rect 1200 1829 1226 1859
rect 1256 1829 1263 1859
rect 1051 1822 1263 1829
rect 1611 1859 1767 1866
rect 1611 1829 1618 1859
rect 1648 1829 1674 1859
rect 1704 1829 1730 1859
rect 1760 1829 1767 1859
rect 1611 1822 1767 1829
rect 2003 1859 2103 1866
rect 2003 1829 2010 1859
rect 2040 1829 2066 1859
rect 2096 1829 2103 1859
rect 2003 1822 2103 1829
rect 2315 1859 2415 1866
rect 2315 1829 2322 1859
rect 2352 1829 2378 1859
rect 2408 1829 2415 1859
rect 2315 1822 2415 1829
rect 2763 1859 2975 1866
rect 2763 1829 2770 1859
rect 2800 1829 2826 1859
rect 2856 1829 2882 1859
rect 2912 1829 2938 1859
rect 2968 1829 2975 1859
rect 2763 1822 2975 1829
rect 3323 1859 3479 1866
rect 3323 1829 3330 1859
rect 3360 1829 3386 1859
rect 3416 1829 3442 1859
rect 3472 1829 3479 1859
rect 3323 1822 3479 1829
rect 3715 1859 3815 1866
rect 3715 1829 3722 1859
rect 3752 1829 3778 1859
rect 3808 1829 3815 1859
rect 3715 1822 3815 1829
rect 4027 1859 4127 1866
rect 4027 1829 4034 1859
rect 4064 1829 4090 1859
rect 4120 1829 4127 1859
rect 4027 1822 4127 1829
rect 4475 1859 4687 1866
rect 4475 1829 4482 1859
rect 4512 1829 4538 1859
rect 4568 1829 4594 1859
rect 4624 1829 4650 1859
rect 4680 1829 4687 1859
rect 4475 1822 4687 1829
rect 5035 1859 5191 1866
rect 5035 1829 5042 1859
rect 5072 1829 5098 1859
rect 5128 1829 5154 1859
rect 5184 1829 5191 1859
rect 5035 1822 5191 1829
rect 5427 1859 5527 1866
rect 5427 1829 5434 1859
rect 5464 1829 5490 1859
rect 5520 1829 5527 1859
rect 5427 1822 5527 1829
rect 5739 1859 5839 1866
rect 5739 1829 5746 1859
rect 5776 1829 5802 1859
rect 5832 1829 5839 1859
rect 5739 1822 5839 1829
rect 6187 1859 6399 1866
rect 6187 1829 6194 1859
rect 6224 1829 6250 1859
rect 6280 1829 6306 1859
rect 6336 1829 6362 1859
rect 6392 1829 6399 1859
rect 6187 1822 6399 1829
rect 6747 1859 6903 1866
rect 6747 1829 6754 1859
rect 6784 1829 6810 1859
rect 6840 1829 6866 1859
rect 6896 1829 6903 1859
rect 6747 1822 6903 1829
rect 7139 1859 7239 1866
rect 7139 1829 7146 1859
rect 7176 1829 7202 1859
rect 7232 1829 7239 1859
rect 7139 1822 7239 1829
rect 7451 1859 7551 1866
rect 7451 1829 7458 1859
rect 7488 1829 7514 1859
rect 7544 1829 7551 1859
rect 7451 1822 7551 1829
rect 7899 1859 8111 1866
rect 7899 1829 7906 1859
rect 7936 1829 7962 1859
rect 7992 1829 8018 1859
rect 8048 1829 8074 1859
rect 8104 1829 8111 1859
rect 7899 1822 8111 1829
rect 8459 1859 8615 1866
rect 8459 1829 8466 1859
rect 8496 1829 8522 1859
rect 8552 1829 8578 1859
rect 8608 1829 8615 1859
rect 8459 1822 8615 1829
rect 8851 1859 8951 1866
rect 8851 1829 8858 1859
rect 8888 1829 8914 1859
rect 8944 1829 8951 1859
rect 8851 1822 8951 1829
rect 9250 1850 9300 2253
rect 9400 2000 9450 2553
rect 9400 1950 10550 2000
rect 9250 1800 10400 1850
rect -150 1185 -100 1800
rect 211 1609 311 1616
rect 211 1579 218 1609
rect 248 1579 274 1609
rect 304 1579 311 1609
rect 211 1572 311 1579
rect 547 1609 703 1616
rect 547 1579 554 1609
rect 584 1579 610 1609
rect 640 1579 666 1609
rect 696 1579 703 1609
rect 547 1572 703 1579
rect 1051 1609 1263 1616
rect 1051 1579 1058 1609
rect 1088 1579 1114 1609
rect 1144 1579 1170 1609
rect 1200 1579 1226 1609
rect 1256 1579 1263 1609
rect 1051 1572 1263 1579
rect 1611 1609 1711 1616
rect 1611 1579 1618 1609
rect 1648 1579 1674 1609
rect 1704 1579 1711 1609
rect 1611 1572 1711 1579
rect 1923 1609 2023 1616
rect 1923 1579 1930 1609
rect 1960 1579 1986 1609
rect 2016 1579 2023 1609
rect 1923 1572 2023 1579
rect 2259 1609 2415 1616
rect 2259 1579 2266 1609
rect 2296 1579 2322 1609
rect 2352 1579 2378 1609
rect 2408 1579 2415 1609
rect 2259 1572 2415 1579
rect 2763 1609 2975 1616
rect 2763 1579 2770 1609
rect 2800 1579 2826 1609
rect 2856 1579 2882 1609
rect 2912 1579 2938 1609
rect 2968 1579 2975 1609
rect 2763 1572 2975 1579
rect 3323 1609 3423 1616
rect 3323 1579 3330 1609
rect 3360 1579 3386 1609
rect 3416 1579 3423 1609
rect 3323 1572 3423 1579
rect 3635 1609 3735 1616
rect 3635 1579 3642 1609
rect 3672 1579 3698 1609
rect 3728 1579 3735 1609
rect 3635 1572 3735 1579
rect 3971 1609 4127 1616
rect 3971 1579 3978 1609
rect 4008 1579 4034 1609
rect 4064 1579 4090 1609
rect 4120 1579 4127 1609
rect 3971 1572 4127 1579
rect 4475 1609 4687 1616
rect 4475 1579 4482 1609
rect 4512 1579 4538 1609
rect 4568 1579 4594 1609
rect 4624 1579 4650 1609
rect 4680 1579 4687 1609
rect 4475 1572 4687 1579
rect 5035 1609 5135 1616
rect 5035 1579 5042 1609
rect 5072 1579 5098 1609
rect 5128 1579 5135 1609
rect 5035 1572 5135 1579
rect 5347 1609 5447 1616
rect 5347 1579 5354 1609
rect 5384 1579 5410 1609
rect 5440 1579 5447 1609
rect 5347 1572 5447 1579
rect 5683 1609 5839 1616
rect 5683 1579 5690 1609
rect 5720 1579 5746 1609
rect 5776 1579 5802 1609
rect 5832 1579 5839 1609
rect 5683 1572 5839 1579
rect 6187 1609 6399 1616
rect 6187 1579 6194 1609
rect 6224 1579 6250 1609
rect 6280 1579 6306 1609
rect 6336 1579 6362 1609
rect 6392 1579 6399 1609
rect 6187 1572 6399 1579
rect 6747 1609 6847 1616
rect 6747 1579 6754 1609
rect 6784 1579 6810 1609
rect 6840 1579 6847 1609
rect 6747 1572 6847 1579
rect 7059 1609 7159 1616
rect 7059 1579 7066 1609
rect 7096 1579 7122 1609
rect 7152 1579 7159 1609
rect 7059 1572 7159 1579
rect 7395 1609 7551 1616
rect 7395 1579 7402 1609
rect 7432 1579 7458 1609
rect 7488 1579 7514 1609
rect 7544 1579 7551 1609
rect 7395 1572 7551 1579
rect 7899 1609 8111 1616
rect 7899 1579 7906 1609
rect 7936 1579 7962 1609
rect 7992 1579 8018 1609
rect 8048 1579 8074 1609
rect 8104 1579 8111 1609
rect 7899 1572 8111 1579
rect 8459 1609 8559 1616
rect 8459 1579 8466 1609
rect 8496 1579 8522 1609
rect 8552 1579 8559 1609
rect 8459 1572 8559 1579
rect 8771 1609 8871 1616
rect 8771 1579 8778 1609
rect 8808 1579 8834 1609
rect 8864 1579 8871 1609
rect 8771 1572 8871 1579
rect 9107 1609 9263 1616
rect 9107 1579 9114 1609
rect 9144 1579 9170 1609
rect 9200 1579 9226 1609
rect 9256 1579 9263 1609
rect 9107 1572 9263 1579
rect 9611 1609 9823 1616
rect 9611 1579 9618 1609
rect 9648 1579 9674 1609
rect 9704 1579 9730 1609
rect 9760 1579 9786 1609
rect 9816 1579 9823 1609
rect 9611 1572 9823 1579
rect 10171 1609 10271 1616
rect 10171 1579 10178 1609
rect 10208 1579 10234 1609
rect 10264 1579 10271 1609
rect 10171 1572 10271 1579
rect 10350 1185 10400 1800
rect -150 1135 0 1185
rect 10200 1135 10400 1185
rect 10500 885 10550 1950
rect -300 835 129 885
rect 10222 835 10550 885
<< via1 >>
rect 610 1829 640 1859
rect 666 1829 696 1859
rect 1058 1829 1088 1859
rect 1114 1829 1144 1859
rect 1170 1829 1200 1859
rect 1226 1829 1256 1859
rect 1618 1829 1648 1859
rect 1674 1829 1704 1859
rect 1730 1829 1760 1859
rect 2010 1829 2040 1859
rect 2066 1829 2096 1859
rect 2322 1829 2352 1859
rect 2378 1829 2408 1859
rect 2770 1829 2800 1859
rect 2826 1829 2856 1859
rect 2882 1829 2912 1859
rect 2938 1829 2968 1859
rect 3330 1829 3360 1859
rect 3386 1829 3416 1859
rect 3442 1829 3472 1859
rect 3722 1829 3752 1859
rect 3778 1829 3808 1859
rect 4034 1829 4064 1859
rect 4090 1829 4120 1859
rect 4482 1829 4512 1859
rect 4538 1829 4568 1859
rect 4594 1829 4624 1859
rect 4650 1829 4680 1859
rect 5042 1829 5072 1859
rect 5098 1829 5128 1859
rect 5154 1829 5184 1859
rect 5434 1829 5464 1859
rect 5490 1829 5520 1859
rect 5746 1829 5776 1859
rect 5802 1829 5832 1859
rect 6194 1829 6224 1859
rect 6250 1829 6280 1859
rect 6306 1829 6336 1859
rect 6362 1829 6392 1859
rect 6754 1829 6784 1859
rect 6810 1829 6840 1859
rect 6866 1829 6896 1859
rect 7146 1829 7176 1859
rect 7202 1829 7232 1859
rect 7458 1829 7488 1859
rect 7514 1829 7544 1859
rect 7906 1829 7936 1859
rect 7962 1829 7992 1859
rect 8018 1829 8048 1859
rect 8074 1829 8104 1859
rect 8466 1829 8496 1859
rect 8522 1829 8552 1859
rect 8578 1829 8608 1859
rect 8858 1829 8888 1859
rect 8914 1829 8944 1859
rect 218 1579 248 1609
rect 274 1579 304 1609
rect 554 1579 584 1609
rect 610 1579 640 1609
rect 666 1579 696 1609
rect 1058 1579 1088 1609
rect 1114 1579 1144 1609
rect 1170 1579 1200 1609
rect 1226 1579 1256 1609
rect 1618 1579 1648 1609
rect 1674 1579 1704 1609
rect 1930 1579 1960 1609
rect 1986 1579 2016 1609
rect 2266 1579 2296 1609
rect 2322 1579 2352 1609
rect 2378 1579 2408 1609
rect 2770 1579 2800 1609
rect 2826 1579 2856 1609
rect 2882 1579 2912 1609
rect 2938 1579 2968 1609
rect 3330 1579 3360 1609
rect 3386 1579 3416 1609
rect 3642 1579 3672 1609
rect 3698 1579 3728 1609
rect 3978 1579 4008 1609
rect 4034 1579 4064 1609
rect 4090 1579 4120 1609
rect 4482 1579 4512 1609
rect 4538 1579 4568 1609
rect 4594 1579 4624 1609
rect 4650 1579 4680 1609
rect 5042 1579 5072 1609
rect 5098 1579 5128 1609
rect 5354 1579 5384 1609
rect 5410 1579 5440 1609
rect 5690 1579 5720 1609
rect 5746 1579 5776 1609
rect 5802 1579 5832 1609
rect 6194 1579 6224 1609
rect 6250 1579 6280 1609
rect 6306 1579 6336 1609
rect 6362 1579 6392 1609
rect 6754 1579 6784 1609
rect 6810 1579 6840 1609
rect 7066 1579 7096 1609
rect 7122 1579 7152 1609
rect 7402 1579 7432 1609
rect 7458 1579 7488 1609
rect 7514 1579 7544 1609
rect 7906 1579 7936 1609
rect 7962 1579 7992 1609
rect 8018 1579 8048 1609
rect 8074 1579 8104 1609
rect 8466 1579 8496 1609
rect 8522 1579 8552 1609
rect 8778 1579 8808 1609
rect 8834 1579 8864 1609
rect 9114 1579 9144 1609
rect 9170 1579 9200 1609
rect 9226 1579 9256 1609
rect 9618 1579 9648 1609
rect 9674 1579 9704 1609
rect 9730 1579 9760 1609
rect 9786 1579 9816 1609
rect 10178 1579 10208 1609
rect 10234 1579 10264 1609
<< metal2 >>
rect 603 1861 703 1866
rect 603 1827 608 1861
rect 642 1827 664 1861
rect 698 1827 703 1861
rect 603 1822 703 1827
rect 1051 1861 1263 1866
rect 1051 1827 1056 1861
rect 1090 1827 1112 1861
rect 1146 1827 1168 1861
rect 1202 1827 1224 1861
rect 1258 1827 1263 1861
rect 1051 1822 1263 1827
rect 1611 1861 1767 1866
rect 1611 1827 1616 1861
rect 1650 1827 1672 1861
rect 1706 1827 1728 1861
rect 1762 1827 1767 1861
rect 1611 1822 1767 1827
rect 2003 1861 2103 1866
rect 2003 1827 2008 1861
rect 2042 1827 2064 1861
rect 2098 1827 2103 1861
rect 2003 1822 2103 1827
rect 2315 1861 2415 1866
rect 2315 1827 2320 1861
rect 2354 1827 2376 1861
rect 2410 1827 2415 1861
rect 2315 1822 2415 1827
rect 2763 1861 2975 1866
rect 2763 1827 2768 1861
rect 2802 1827 2824 1861
rect 2858 1827 2880 1861
rect 2914 1827 2936 1861
rect 2970 1827 2975 1861
rect 2763 1822 2975 1827
rect 3323 1861 3479 1866
rect 3323 1827 3328 1861
rect 3362 1827 3384 1861
rect 3418 1827 3440 1861
rect 3474 1827 3479 1861
rect 3323 1822 3479 1827
rect 3715 1861 3815 1866
rect 3715 1827 3720 1861
rect 3754 1827 3776 1861
rect 3810 1827 3815 1861
rect 3715 1822 3815 1827
rect 4027 1861 4127 1866
rect 4027 1827 4032 1861
rect 4066 1827 4088 1861
rect 4122 1827 4127 1861
rect 4027 1822 4127 1827
rect 4475 1861 4687 1866
rect 4475 1827 4480 1861
rect 4514 1827 4536 1861
rect 4570 1827 4592 1861
rect 4626 1827 4648 1861
rect 4682 1827 4687 1861
rect 4475 1822 4687 1827
rect 5035 1861 5191 1866
rect 5035 1827 5040 1861
rect 5074 1827 5096 1861
rect 5130 1827 5152 1861
rect 5186 1827 5191 1861
rect 5035 1822 5191 1827
rect 5427 1861 5527 1866
rect 5427 1827 5432 1861
rect 5466 1827 5488 1861
rect 5522 1827 5527 1861
rect 5427 1822 5527 1827
rect 5739 1861 5839 1866
rect 5739 1827 5744 1861
rect 5778 1827 5800 1861
rect 5834 1827 5839 1861
rect 5739 1822 5839 1827
rect 6187 1861 6399 1866
rect 6187 1827 6192 1861
rect 6226 1827 6248 1861
rect 6282 1827 6304 1861
rect 6338 1827 6360 1861
rect 6394 1827 6399 1861
rect 6187 1822 6399 1827
rect 6747 1861 6903 1866
rect 6747 1827 6752 1861
rect 6786 1827 6808 1861
rect 6842 1827 6864 1861
rect 6898 1827 6903 1861
rect 6747 1822 6903 1827
rect 7139 1861 7239 1866
rect 7139 1827 7144 1861
rect 7178 1827 7200 1861
rect 7234 1827 7239 1861
rect 7139 1822 7239 1827
rect 7451 1861 7551 1866
rect 7451 1827 7456 1861
rect 7490 1827 7512 1861
rect 7546 1827 7551 1861
rect 7451 1822 7551 1827
rect 7899 1861 8111 1866
rect 7899 1827 7904 1861
rect 7938 1827 7960 1861
rect 7994 1827 8016 1861
rect 8050 1827 8072 1861
rect 8106 1827 8111 1861
rect 7899 1822 8111 1827
rect 8459 1861 8615 1866
rect 8459 1827 8464 1861
rect 8498 1827 8520 1861
rect 8554 1827 8576 1861
rect 8610 1827 8615 1861
rect 8459 1822 8615 1827
rect 8851 1861 8951 1866
rect 8851 1827 8856 1861
rect 8890 1827 8912 1861
rect 8946 1827 8951 1861
rect 8851 1822 8951 1827
rect 211 1611 311 1616
rect 211 1577 216 1611
rect 250 1577 272 1611
rect 306 1577 311 1611
rect 211 1572 311 1577
rect 547 1611 703 1616
rect 547 1577 552 1611
rect 586 1577 608 1611
rect 642 1577 664 1611
rect 698 1577 703 1611
rect 547 1572 703 1577
rect 1051 1611 1263 1616
rect 1051 1577 1056 1611
rect 1090 1577 1112 1611
rect 1146 1577 1168 1611
rect 1202 1577 1224 1611
rect 1258 1577 1263 1611
rect 1051 1572 1263 1577
rect 1611 1611 1711 1616
rect 1611 1577 1616 1611
rect 1650 1577 1672 1611
rect 1706 1577 1711 1611
rect 1611 1572 1711 1577
rect 1923 1611 2023 1616
rect 1923 1577 1928 1611
rect 1962 1577 1984 1611
rect 2018 1577 2023 1611
rect 1923 1572 2023 1577
rect 2259 1611 2415 1616
rect 2259 1577 2264 1611
rect 2298 1577 2320 1611
rect 2354 1577 2376 1611
rect 2410 1577 2415 1611
rect 2259 1572 2415 1577
rect 2763 1611 2975 1616
rect 2763 1577 2768 1611
rect 2802 1577 2824 1611
rect 2858 1577 2880 1611
rect 2914 1577 2936 1611
rect 2970 1577 2975 1611
rect 2763 1572 2975 1577
rect 3323 1611 3423 1616
rect 3323 1577 3328 1611
rect 3362 1577 3384 1611
rect 3418 1577 3423 1611
rect 3323 1572 3423 1577
rect 3635 1611 3735 1616
rect 3635 1577 3640 1611
rect 3674 1577 3696 1611
rect 3730 1577 3735 1611
rect 3635 1572 3735 1577
rect 3971 1611 4127 1616
rect 3971 1577 3976 1611
rect 4010 1577 4032 1611
rect 4066 1577 4088 1611
rect 4122 1577 4127 1611
rect 3971 1572 4127 1577
rect 4475 1611 4687 1616
rect 4475 1577 4480 1611
rect 4514 1577 4536 1611
rect 4570 1577 4592 1611
rect 4626 1577 4648 1611
rect 4682 1577 4687 1611
rect 4475 1572 4687 1577
rect 5035 1611 5135 1616
rect 5035 1577 5040 1611
rect 5074 1577 5096 1611
rect 5130 1577 5135 1611
rect 5035 1572 5135 1577
rect 5347 1611 5447 1616
rect 5347 1577 5352 1611
rect 5386 1577 5408 1611
rect 5442 1577 5447 1611
rect 5347 1572 5447 1577
rect 5683 1611 5839 1616
rect 5683 1577 5688 1611
rect 5722 1577 5744 1611
rect 5778 1577 5800 1611
rect 5834 1577 5839 1611
rect 5683 1572 5839 1577
rect 6187 1611 6399 1616
rect 6187 1577 6192 1611
rect 6226 1577 6248 1611
rect 6282 1577 6304 1611
rect 6338 1577 6360 1611
rect 6394 1577 6399 1611
rect 6187 1572 6399 1577
rect 6747 1611 6847 1616
rect 6747 1577 6752 1611
rect 6786 1577 6808 1611
rect 6842 1577 6847 1611
rect 6747 1572 6847 1577
rect 7059 1611 7159 1616
rect 7059 1577 7064 1611
rect 7098 1577 7120 1611
rect 7154 1577 7159 1611
rect 7059 1572 7159 1577
rect 7395 1611 7551 1616
rect 7395 1577 7400 1611
rect 7434 1577 7456 1611
rect 7490 1577 7512 1611
rect 7546 1577 7551 1611
rect 7395 1572 7551 1577
rect 7899 1611 8111 1616
rect 7899 1577 7904 1611
rect 7938 1577 7960 1611
rect 7994 1577 8016 1611
rect 8050 1577 8072 1611
rect 8106 1577 8111 1611
rect 7899 1572 8111 1577
rect 8459 1611 8559 1616
rect 8459 1577 8464 1611
rect 8498 1577 8520 1611
rect 8554 1577 8559 1611
rect 8459 1572 8559 1577
rect 8771 1611 8871 1616
rect 8771 1577 8776 1611
rect 8810 1577 8832 1611
rect 8866 1577 8871 1611
rect 8771 1572 8871 1577
rect 9107 1611 9263 1616
rect 9107 1577 9112 1611
rect 9146 1577 9168 1611
rect 9202 1577 9224 1611
rect 9258 1577 9263 1611
rect 9107 1572 9263 1577
rect 9611 1611 9823 1616
rect 9611 1577 9616 1611
rect 9650 1577 9672 1611
rect 9706 1577 9728 1611
rect 9762 1577 9784 1611
rect 9818 1577 9823 1611
rect 9611 1572 9823 1577
rect 10171 1611 10271 1616
rect 10171 1577 10176 1611
rect 10210 1577 10232 1611
rect 10266 1577 10271 1611
rect 10171 1572 10271 1577
<< via2 >>
rect 608 1859 642 1861
rect 608 1829 610 1859
rect 610 1829 640 1859
rect 640 1829 642 1859
rect 608 1827 642 1829
rect 664 1859 698 1861
rect 664 1829 666 1859
rect 666 1829 696 1859
rect 696 1829 698 1859
rect 664 1827 698 1829
rect 1056 1859 1090 1861
rect 1056 1829 1058 1859
rect 1058 1829 1088 1859
rect 1088 1829 1090 1859
rect 1056 1827 1090 1829
rect 1112 1859 1146 1861
rect 1112 1829 1114 1859
rect 1114 1829 1144 1859
rect 1144 1829 1146 1859
rect 1112 1827 1146 1829
rect 1168 1859 1202 1861
rect 1168 1829 1170 1859
rect 1170 1829 1200 1859
rect 1200 1829 1202 1859
rect 1168 1827 1202 1829
rect 1224 1859 1258 1861
rect 1224 1829 1226 1859
rect 1226 1829 1256 1859
rect 1256 1829 1258 1859
rect 1224 1827 1258 1829
rect 1616 1859 1650 1861
rect 1616 1829 1618 1859
rect 1618 1829 1648 1859
rect 1648 1829 1650 1859
rect 1616 1827 1650 1829
rect 1672 1859 1706 1861
rect 1672 1829 1674 1859
rect 1674 1829 1704 1859
rect 1704 1829 1706 1859
rect 1672 1827 1706 1829
rect 1728 1859 1762 1861
rect 1728 1829 1730 1859
rect 1730 1829 1760 1859
rect 1760 1829 1762 1859
rect 1728 1827 1762 1829
rect 2008 1859 2042 1861
rect 2008 1829 2010 1859
rect 2010 1829 2040 1859
rect 2040 1829 2042 1859
rect 2008 1827 2042 1829
rect 2064 1859 2098 1861
rect 2064 1829 2066 1859
rect 2066 1829 2096 1859
rect 2096 1829 2098 1859
rect 2064 1827 2098 1829
rect 2320 1859 2354 1861
rect 2320 1829 2322 1859
rect 2322 1829 2352 1859
rect 2352 1829 2354 1859
rect 2320 1827 2354 1829
rect 2376 1859 2410 1861
rect 2376 1829 2378 1859
rect 2378 1829 2408 1859
rect 2408 1829 2410 1859
rect 2376 1827 2410 1829
rect 2768 1859 2802 1861
rect 2768 1829 2770 1859
rect 2770 1829 2800 1859
rect 2800 1829 2802 1859
rect 2768 1827 2802 1829
rect 2824 1859 2858 1861
rect 2824 1829 2826 1859
rect 2826 1829 2856 1859
rect 2856 1829 2858 1859
rect 2824 1827 2858 1829
rect 2880 1859 2914 1861
rect 2880 1829 2882 1859
rect 2882 1829 2912 1859
rect 2912 1829 2914 1859
rect 2880 1827 2914 1829
rect 2936 1859 2970 1861
rect 2936 1829 2938 1859
rect 2938 1829 2968 1859
rect 2968 1829 2970 1859
rect 2936 1827 2970 1829
rect 3328 1859 3362 1861
rect 3328 1829 3330 1859
rect 3330 1829 3360 1859
rect 3360 1829 3362 1859
rect 3328 1827 3362 1829
rect 3384 1859 3418 1861
rect 3384 1829 3386 1859
rect 3386 1829 3416 1859
rect 3416 1829 3418 1859
rect 3384 1827 3418 1829
rect 3440 1859 3474 1861
rect 3440 1829 3442 1859
rect 3442 1829 3472 1859
rect 3472 1829 3474 1859
rect 3440 1827 3474 1829
rect 3720 1859 3754 1861
rect 3720 1829 3722 1859
rect 3722 1829 3752 1859
rect 3752 1829 3754 1859
rect 3720 1827 3754 1829
rect 3776 1859 3810 1861
rect 3776 1829 3778 1859
rect 3778 1829 3808 1859
rect 3808 1829 3810 1859
rect 3776 1827 3810 1829
rect 4032 1859 4066 1861
rect 4032 1829 4034 1859
rect 4034 1829 4064 1859
rect 4064 1829 4066 1859
rect 4032 1827 4066 1829
rect 4088 1859 4122 1861
rect 4088 1829 4090 1859
rect 4090 1829 4120 1859
rect 4120 1829 4122 1859
rect 4088 1827 4122 1829
rect 4480 1859 4514 1861
rect 4480 1829 4482 1859
rect 4482 1829 4512 1859
rect 4512 1829 4514 1859
rect 4480 1827 4514 1829
rect 4536 1859 4570 1861
rect 4536 1829 4538 1859
rect 4538 1829 4568 1859
rect 4568 1829 4570 1859
rect 4536 1827 4570 1829
rect 4592 1859 4626 1861
rect 4592 1829 4594 1859
rect 4594 1829 4624 1859
rect 4624 1829 4626 1859
rect 4592 1827 4626 1829
rect 4648 1859 4682 1861
rect 4648 1829 4650 1859
rect 4650 1829 4680 1859
rect 4680 1829 4682 1859
rect 4648 1827 4682 1829
rect 5040 1859 5074 1861
rect 5040 1829 5042 1859
rect 5042 1829 5072 1859
rect 5072 1829 5074 1859
rect 5040 1827 5074 1829
rect 5096 1859 5130 1861
rect 5096 1829 5098 1859
rect 5098 1829 5128 1859
rect 5128 1829 5130 1859
rect 5096 1827 5130 1829
rect 5152 1859 5186 1861
rect 5152 1829 5154 1859
rect 5154 1829 5184 1859
rect 5184 1829 5186 1859
rect 5152 1827 5186 1829
rect 5432 1859 5466 1861
rect 5432 1829 5434 1859
rect 5434 1829 5464 1859
rect 5464 1829 5466 1859
rect 5432 1827 5466 1829
rect 5488 1859 5522 1861
rect 5488 1829 5490 1859
rect 5490 1829 5520 1859
rect 5520 1829 5522 1859
rect 5488 1827 5522 1829
rect 5744 1859 5778 1861
rect 5744 1829 5746 1859
rect 5746 1829 5776 1859
rect 5776 1829 5778 1859
rect 5744 1827 5778 1829
rect 5800 1859 5834 1861
rect 5800 1829 5802 1859
rect 5802 1829 5832 1859
rect 5832 1829 5834 1859
rect 5800 1827 5834 1829
rect 6192 1859 6226 1861
rect 6192 1829 6194 1859
rect 6194 1829 6224 1859
rect 6224 1829 6226 1859
rect 6192 1827 6226 1829
rect 6248 1859 6282 1861
rect 6248 1829 6250 1859
rect 6250 1829 6280 1859
rect 6280 1829 6282 1859
rect 6248 1827 6282 1829
rect 6304 1859 6338 1861
rect 6304 1829 6306 1859
rect 6306 1829 6336 1859
rect 6336 1829 6338 1859
rect 6304 1827 6338 1829
rect 6360 1859 6394 1861
rect 6360 1829 6362 1859
rect 6362 1829 6392 1859
rect 6392 1829 6394 1859
rect 6360 1827 6394 1829
rect 6752 1859 6786 1861
rect 6752 1829 6754 1859
rect 6754 1829 6784 1859
rect 6784 1829 6786 1859
rect 6752 1827 6786 1829
rect 6808 1859 6842 1861
rect 6808 1829 6810 1859
rect 6810 1829 6840 1859
rect 6840 1829 6842 1859
rect 6808 1827 6842 1829
rect 6864 1859 6898 1861
rect 6864 1829 6866 1859
rect 6866 1829 6896 1859
rect 6896 1829 6898 1859
rect 6864 1827 6898 1829
rect 7144 1859 7178 1861
rect 7144 1829 7146 1859
rect 7146 1829 7176 1859
rect 7176 1829 7178 1859
rect 7144 1827 7178 1829
rect 7200 1859 7234 1861
rect 7200 1829 7202 1859
rect 7202 1829 7232 1859
rect 7232 1829 7234 1859
rect 7200 1827 7234 1829
rect 7456 1859 7490 1861
rect 7456 1829 7458 1859
rect 7458 1829 7488 1859
rect 7488 1829 7490 1859
rect 7456 1827 7490 1829
rect 7512 1859 7546 1861
rect 7512 1829 7514 1859
rect 7514 1829 7544 1859
rect 7544 1829 7546 1859
rect 7512 1827 7546 1829
rect 7904 1859 7938 1861
rect 7904 1829 7906 1859
rect 7906 1829 7936 1859
rect 7936 1829 7938 1859
rect 7904 1827 7938 1829
rect 7960 1859 7994 1861
rect 7960 1829 7962 1859
rect 7962 1829 7992 1859
rect 7992 1829 7994 1859
rect 7960 1827 7994 1829
rect 8016 1859 8050 1861
rect 8016 1829 8018 1859
rect 8018 1829 8048 1859
rect 8048 1829 8050 1859
rect 8016 1827 8050 1829
rect 8072 1859 8106 1861
rect 8072 1829 8074 1859
rect 8074 1829 8104 1859
rect 8104 1829 8106 1859
rect 8072 1827 8106 1829
rect 8464 1859 8498 1861
rect 8464 1829 8466 1859
rect 8466 1829 8496 1859
rect 8496 1829 8498 1859
rect 8464 1827 8498 1829
rect 8520 1859 8554 1861
rect 8520 1829 8522 1859
rect 8522 1829 8552 1859
rect 8552 1829 8554 1859
rect 8520 1827 8554 1829
rect 8576 1859 8610 1861
rect 8576 1829 8578 1859
rect 8578 1829 8608 1859
rect 8608 1829 8610 1859
rect 8576 1827 8610 1829
rect 8856 1859 8890 1861
rect 8856 1829 8858 1859
rect 8858 1829 8888 1859
rect 8888 1829 8890 1859
rect 8856 1827 8890 1829
rect 8912 1859 8946 1861
rect 8912 1829 8914 1859
rect 8914 1829 8944 1859
rect 8944 1829 8946 1859
rect 8912 1827 8946 1829
rect 216 1609 250 1611
rect 216 1579 218 1609
rect 218 1579 248 1609
rect 248 1579 250 1609
rect 216 1577 250 1579
rect 272 1609 306 1611
rect 272 1579 274 1609
rect 274 1579 304 1609
rect 304 1579 306 1609
rect 272 1577 306 1579
rect 552 1609 586 1611
rect 552 1579 554 1609
rect 554 1579 584 1609
rect 584 1579 586 1609
rect 552 1577 586 1579
rect 608 1609 642 1611
rect 608 1579 610 1609
rect 610 1579 640 1609
rect 640 1579 642 1609
rect 608 1577 642 1579
rect 664 1609 698 1611
rect 664 1579 666 1609
rect 666 1579 696 1609
rect 696 1579 698 1609
rect 664 1577 698 1579
rect 1056 1609 1090 1611
rect 1056 1579 1058 1609
rect 1058 1579 1088 1609
rect 1088 1579 1090 1609
rect 1056 1577 1090 1579
rect 1112 1609 1146 1611
rect 1112 1579 1114 1609
rect 1114 1579 1144 1609
rect 1144 1579 1146 1609
rect 1112 1577 1146 1579
rect 1168 1609 1202 1611
rect 1168 1579 1170 1609
rect 1170 1579 1200 1609
rect 1200 1579 1202 1609
rect 1168 1577 1202 1579
rect 1224 1609 1258 1611
rect 1224 1579 1226 1609
rect 1226 1579 1256 1609
rect 1256 1579 1258 1609
rect 1224 1577 1258 1579
rect 1616 1609 1650 1611
rect 1616 1579 1618 1609
rect 1618 1579 1648 1609
rect 1648 1579 1650 1609
rect 1616 1577 1650 1579
rect 1672 1609 1706 1611
rect 1672 1579 1674 1609
rect 1674 1579 1704 1609
rect 1704 1579 1706 1609
rect 1672 1577 1706 1579
rect 1928 1609 1962 1611
rect 1928 1579 1930 1609
rect 1930 1579 1960 1609
rect 1960 1579 1962 1609
rect 1928 1577 1962 1579
rect 1984 1609 2018 1611
rect 1984 1579 1986 1609
rect 1986 1579 2016 1609
rect 2016 1579 2018 1609
rect 1984 1577 2018 1579
rect 2264 1609 2298 1611
rect 2264 1579 2266 1609
rect 2266 1579 2296 1609
rect 2296 1579 2298 1609
rect 2264 1577 2298 1579
rect 2320 1609 2354 1611
rect 2320 1579 2322 1609
rect 2322 1579 2352 1609
rect 2352 1579 2354 1609
rect 2320 1577 2354 1579
rect 2376 1609 2410 1611
rect 2376 1579 2378 1609
rect 2378 1579 2408 1609
rect 2408 1579 2410 1609
rect 2376 1577 2410 1579
rect 2768 1609 2802 1611
rect 2768 1579 2770 1609
rect 2770 1579 2800 1609
rect 2800 1579 2802 1609
rect 2768 1577 2802 1579
rect 2824 1609 2858 1611
rect 2824 1579 2826 1609
rect 2826 1579 2856 1609
rect 2856 1579 2858 1609
rect 2824 1577 2858 1579
rect 2880 1609 2914 1611
rect 2880 1579 2882 1609
rect 2882 1579 2912 1609
rect 2912 1579 2914 1609
rect 2880 1577 2914 1579
rect 2936 1609 2970 1611
rect 2936 1579 2938 1609
rect 2938 1579 2968 1609
rect 2968 1579 2970 1609
rect 2936 1577 2970 1579
rect 3328 1609 3362 1611
rect 3328 1579 3330 1609
rect 3330 1579 3360 1609
rect 3360 1579 3362 1609
rect 3328 1577 3362 1579
rect 3384 1609 3418 1611
rect 3384 1579 3386 1609
rect 3386 1579 3416 1609
rect 3416 1579 3418 1609
rect 3384 1577 3418 1579
rect 3640 1609 3674 1611
rect 3640 1579 3642 1609
rect 3642 1579 3672 1609
rect 3672 1579 3674 1609
rect 3640 1577 3674 1579
rect 3696 1609 3730 1611
rect 3696 1579 3698 1609
rect 3698 1579 3728 1609
rect 3728 1579 3730 1609
rect 3696 1577 3730 1579
rect 3976 1609 4010 1611
rect 3976 1579 3978 1609
rect 3978 1579 4008 1609
rect 4008 1579 4010 1609
rect 3976 1577 4010 1579
rect 4032 1609 4066 1611
rect 4032 1579 4034 1609
rect 4034 1579 4064 1609
rect 4064 1579 4066 1609
rect 4032 1577 4066 1579
rect 4088 1609 4122 1611
rect 4088 1579 4090 1609
rect 4090 1579 4120 1609
rect 4120 1579 4122 1609
rect 4088 1577 4122 1579
rect 4480 1609 4514 1611
rect 4480 1579 4482 1609
rect 4482 1579 4512 1609
rect 4512 1579 4514 1609
rect 4480 1577 4514 1579
rect 4536 1609 4570 1611
rect 4536 1579 4538 1609
rect 4538 1579 4568 1609
rect 4568 1579 4570 1609
rect 4536 1577 4570 1579
rect 4592 1609 4626 1611
rect 4592 1579 4594 1609
rect 4594 1579 4624 1609
rect 4624 1579 4626 1609
rect 4592 1577 4626 1579
rect 4648 1609 4682 1611
rect 4648 1579 4650 1609
rect 4650 1579 4680 1609
rect 4680 1579 4682 1609
rect 4648 1577 4682 1579
rect 5040 1609 5074 1611
rect 5040 1579 5042 1609
rect 5042 1579 5072 1609
rect 5072 1579 5074 1609
rect 5040 1577 5074 1579
rect 5096 1609 5130 1611
rect 5096 1579 5098 1609
rect 5098 1579 5128 1609
rect 5128 1579 5130 1609
rect 5096 1577 5130 1579
rect 5352 1609 5386 1611
rect 5352 1579 5354 1609
rect 5354 1579 5384 1609
rect 5384 1579 5386 1609
rect 5352 1577 5386 1579
rect 5408 1609 5442 1611
rect 5408 1579 5410 1609
rect 5410 1579 5440 1609
rect 5440 1579 5442 1609
rect 5408 1577 5442 1579
rect 5688 1609 5722 1611
rect 5688 1579 5690 1609
rect 5690 1579 5720 1609
rect 5720 1579 5722 1609
rect 5688 1577 5722 1579
rect 5744 1609 5778 1611
rect 5744 1579 5746 1609
rect 5746 1579 5776 1609
rect 5776 1579 5778 1609
rect 5744 1577 5778 1579
rect 5800 1609 5834 1611
rect 5800 1579 5802 1609
rect 5802 1579 5832 1609
rect 5832 1579 5834 1609
rect 5800 1577 5834 1579
rect 6192 1609 6226 1611
rect 6192 1579 6194 1609
rect 6194 1579 6224 1609
rect 6224 1579 6226 1609
rect 6192 1577 6226 1579
rect 6248 1609 6282 1611
rect 6248 1579 6250 1609
rect 6250 1579 6280 1609
rect 6280 1579 6282 1609
rect 6248 1577 6282 1579
rect 6304 1609 6338 1611
rect 6304 1579 6306 1609
rect 6306 1579 6336 1609
rect 6336 1579 6338 1609
rect 6304 1577 6338 1579
rect 6360 1609 6394 1611
rect 6360 1579 6362 1609
rect 6362 1579 6392 1609
rect 6392 1579 6394 1609
rect 6360 1577 6394 1579
rect 6752 1609 6786 1611
rect 6752 1579 6754 1609
rect 6754 1579 6784 1609
rect 6784 1579 6786 1609
rect 6752 1577 6786 1579
rect 6808 1609 6842 1611
rect 6808 1579 6810 1609
rect 6810 1579 6840 1609
rect 6840 1579 6842 1609
rect 6808 1577 6842 1579
rect 7064 1609 7098 1611
rect 7064 1579 7066 1609
rect 7066 1579 7096 1609
rect 7096 1579 7098 1609
rect 7064 1577 7098 1579
rect 7120 1609 7154 1611
rect 7120 1579 7122 1609
rect 7122 1579 7152 1609
rect 7152 1579 7154 1609
rect 7120 1577 7154 1579
rect 7400 1609 7434 1611
rect 7400 1579 7402 1609
rect 7402 1579 7432 1609
rect 7432 1579 7434 1609
rect 7400 1577 7434 1579
rect 7456 1609 7490 1611
rect 7456 1579 7458 1609
rect 7458 1579 7488 1609
rect 7488 1579 7490 1609
rect 7456 1577 7490 1579
rect 7512 1609 7546 1611
rect 7512 1579 7514 1609
rect 7514 1579 7544 1609
rect 7544 1579 7546 1609
rect 7512 1577 7546 1579
rect 7904 1609 7938 1611
rect 7904 1579 7906 1609
rect 7906 1579 7936 1609
rect 7936 1579 7938 1609
rect 7904 1577 7938 1579
rect 7960 1609 7994 1611
rect 7960 1579 7962 1609
rect 7962 1579 7992 1609
rect 7992 1579 7994 1609
rect 7960 1577 7994 1579
rect 8016 1609 8050 1611
rect 8016 1579 8018 1609
rect 8018 1579 8048 1609
rect 8048 1579 8050 1609
rect 8016 1577 8050 1579
rect 8072 1609 8106 1611
rect 8072 1579 8074 1609
rect 8074 1579 8104 1609
rect 8104 1579 8106 1609
rect 8072 1577 8106 1579
rect 8464 1609 8498 1611
rect 8464 1579 8466 1609
rect 8466 1579 8496 1609
rect 8496 1579 8498 1609
rect 8464 1577 8498 1579
rect 8520 1609 8554 1611
rect 8520 1579 8522 1609
rect 8522 1579 8552 1609
rect 8552 1579 8554 1609
rect 8520 1577 8554 1579
rect 8776 1609 8810 1611
rect 8776 1579 8778 1609
rect 8778 1579 8808 1609
rect 8808 1579 8810 1609
rect 8776 1577 8810 1579
rect 8832 1609 8866 1611
rect 8832 1579 8834 1609
rect 8834 1579 8864 1609
rect 8864 1579 8866 1609
rect 8832 1577 8866 1579
rect 9112 1609 9146 1611
rect 9112 1579 9114 1609
rect 9114 1579 9144 1609
rect 9144 1579 9146 1609
rect 9112 1577 9146 1579
rect 9168 1609 9202 1611
rect 9168 1579 9170 1609
rect 9170 1579 9200 1609
rect 9200 1579 9202 1609
rect 9168 1577 9202 1579
rect 9224 1609 9258 1611
rect 9224 1579 9226 1609
rect 9226 1579 9256 1609
rect 9256 1579 9258 1609
rect 9224 1577 9258 1579
rect 9616 1609 9650 1611
rect 9616 1579 9618 1609
rect 9618 1579 9648 1609
rect 9648 1579 9650 1609
rect 9616 1577 9650 1579
rect 9672 1609 9706 1611
rect 9672 1579 9674 1609
rect 9674 1579 9704 1609
rect 9704 1579 9706 1609
rect 9672 1577 9706 1579
rect 9728 1609 9762 1611
rect 9728 1579 9730 1609
rect 9730 1579 9760 1609
rect 9760 1579 9762 1609
rect 9728 1577 9762 1579
rect 9784 1609 9818 1611
rect 9784 1579 9786 1609
rect 9786 1579 9816 1609
rect 9816 1579 9818 1609
rect 9784 1577 9818 1579
rect 10176 1609 10210 1611
rect 10176 1579 10178 1609
rect 10178 1579 10208 1609
rect 10208 1579 10210 1609
rect 10176 1577 10210 1579
rect 10232 1609 10266 1611
rect 10232 1579 10234 1609
rect 10234 1579 10264 1609
rect 10264 1579 10266 1609
rect 10232 1577 10266 1579
<< metal3 >>
rect 603 1861 703 1866
rect 603 1827 608 1861
rect 642 1827 664 1861
rect 698 1827 703 1861
rect 603 1819 703 1827
rect 1051 1861 1263 1866
rect 1051 1827 1056 1861
rect 1090 1827 1112 1861
rect 1146 1827 1168 1861
rect 1202 1827 1224 1861
rect 1258 1827 1263 1861
rect 1051 1819 1263 1827
rect 1611 1861 1767 1866
rect 1611 1827 1616 1861
rect 1650 1827 1672 1861
rect 1706 1827 1728 1861
rect 1762 1827 1767 1861
rect 1611 1819 1767 1827
rect 2003 1861 2103 1866
rect 2003 1827 2008 1861
rect 2042 1827 2064 1861
rect 2098 1827 2103 1861
rect 2003 1819 2103 1827
rect 2315 1861 2415 1866
rect 2315 1827 2320 1861
rect 2354 1827 2376 1861
rect 2410 1827 2415 1861
rect 2315 1819 2415 1827
rect 2763 1861 2975 1866
rect 2763 1827 2768 1861
rect 2802 1827 2824 1861
rect 2858 1827 2880 1861
rect 2914 1827 2936 1861
rect 2970 1827 2975 1861
rect 2763 1819 2975 1827
rect 3323 1861 3479 1866
rect 3323 1827 3328 1861
rect 3362 1827 3384 1861
rect 3418 1827 3440 1861
rect 3474 1827 3479 1861
rect 3323 1819 3479 1827
rect 3715 1861 3815 1866
rect 3715 1827 3720 1861
rect 3754 1827 3776 1861
rect 3810 1827 3815 1861
rect 3715 1819 3815 1827
rect 4027 1861 4127 1866
rect 4027 1827 4032 1861
rect 4066 1827 4088 1861
rect 4122 1827 4127 1861
rect 4027 1819 4127 1827
rect 4475 1861 4687 1866
rect 4475 1827 4480 1861
rect 4514 1827 4536 1861
rect 4570 1827 4592 1861
rect 4626 1827 4648 1861
rect 4682 1827 4687 1861
rect 4475 1819 4687 1827
rect 5035 1861 5191 1866
rect 5035 1827 5040 1861
rect 5074 1827 5096 1861
rect 5130 1827 5152 1861
rect 5186 1827 5191 1861
rect 5035 1819 5191 1827
rect 5427 1861 5527 1866
rect 5427 1827 5432 1861
rect 5466 1827 5488 1861
rect 5522 1827 5527 1861
rect 5427 1819 5527 1827
rect 5739 1861 5839 1866
rect 5739 1827 5744 1861
rect 5778 1827 5800 1861
rect 5834 1827 5839 1861
rect 5739 1819 5839 1827
rect 6187 1861 6399 1866
rect 6187 1827 6192 1861
rect 6226 1827 6248 1861
rect 6282 1827 6304 1861
rect 6338 1827 6360 1861
rect 6394 1827 6399 1861
rect 6187 1819 6399 1827
rect 6747 1861 6903 1866
rect 6747 1827 6752 1861
rect 6786 1827 6808 1861
rect 6842 1827 6864 1861
rect 6898 1827 6903 1861
rect 6747 1819 6903 1827
rect 7139 1861 7239 1866
rect 7139 1827 7144 1861
rect 7178 1827 7200 1861
rect 7234 1827 7239 1861
rect 7139 1819 7239 1827
rect 7451 1861 7551 1866
rect 7451 1827 7456 1861
rect 7490 1827 7512 1861
rect 7546 1827 7551 1861
rect 7451 1819 7551 1827
rect 7899 1861 8111 1866
rect 7899 1827 7904 1861
rect 7938 1827 7960 1861
rect 7994 1827 8016 1861
rect 8050 1827 8072 1861
rect 8106 1827 8111 1861
rect 7899 1819 8111 1827
rect 8459 1861 8615 1866
rect 8459 1827 8464 1861
rect 8498 1827 8520 1861
rect 8554 1827 8576 1861
rect 8610 1827 8615 1861
rect 8459 1819 8615 1827
rect 8851 1861 8951 1866
rect 8851 1827 8856 1861
rect 8890 1827 8912 1861
rect 8946 1827 8951 1861
rect 8851 1819 8951 1827
rect 0 1619 10272 1819
rect 211 1611 311 1619
rect 211 1577 216 1611
rect 250 1577 272 1611
rect 306 1577 311 1611
rect 211 1572 311 1577
rect 547 1611 703 1619
rect 547 1577 552 1611
rect 586 1577 608 1611
rect 642 1577 664 1611
rect 698 1577 703 1611
rect 547 1572 703 1577
rect 1051 1611 1263 1619
rect 1051 1577 1056 1611
rect 1090 1577 1112 1611
rect 1146 1577 1168 1611
rect 1202 1577 1224 1611
rect 1258 1577 1263 1611
rect 1051 1572 1263 1577
rect 1611 1611 1711 1619
rect 1611 1577 1616 1611
rect 1650 1577 1672 1611
rect 1706 1577 1711 1611
rect 1611 1572 1711 1577
rect 1923 1611 2023 1619
rect 1923 1577 1928 1611
rect 1962 1577 1984 1611
rect 2018 1577 2023 1611
rect 1923 1572 2023 1577
rect 2259 1611 2415 1619
rect 2259 1577 2264 1611
rect 2298 1577 2320 1611
rect 2354 1577 2376 1611
rect 2410 1577 2415 1611
rect 2259 1572 2415 1577
rect 2763 1611 2975 1619
rect 2763 1577 2768 1611
rect 2802 1577 2824 1611
rect 2858 1577 2880 1611
rect 2914 1577 2936 1611
rect 2970 1577 2975 1611
rect 2763 1572 2975 1577
rect 3323 1611 3423 1619
rect 3323 1577 3328 1611
rect 3362 1577 3384 1611
rect 3418 1577 3423 1611
rect 3323 1572 3423 1577
rect 3635 1611 3735 1619
rect 3635 1577 3640 1611
rect 3674 1577 3696 1611
rect 3730 1577 3735 1611
rect 3635 1572 3735 1577
rect 3971 1611 4127 1619
rect 3971 1577 3976 1611
rect 4010 1577 4032 1611
rect 4066 1577 4088 1611
rect 4122 1577 4127 1611
rect 3971 1572 4127 1577
rect 4475 1611 4687 1619
rect 4475 1577 4480 1611
rect 4514 1577 4536 1611
rect 4570 1577 4592 1611
rect 4626 1577 4648 1611
rect 4682 1577 4687 1611
rect 4475 1572 4687 1577
rect 5035 1611 5135 1619
rect 5035 1577 5040 1611
rect 5074 1577 5096 1611
rect 5130 1577 5135 1611
rect 5035 1572 5135 1577
rect 5347 1611 5447 1619
rect 5347 1577 5352 1611
rect 5386 1577 5408 1611
rect 5442 1577 5447 1611
rect 5347 1572 5447 1577
rect 5683 1611 5839 1619
rect 5683 1577 5688 1611
rect 5722 1577 5744 1611
rect 5778 1577 5800 1611
rect 5834 1577 5839 1611
rect 5683 1572 5839 1577
rect 6187 1611 6399 1619
rect 6187 1577 6192 1611
rect 6226 1577 6248 1611
rect 6282 1577 6304 1611
rect 6338 1577 6360 1611
rect 6394 1577 6399 1611
rect 6187 1572 6399 1577
rect 6747 1611 6847 1619
rect 6747 1577 6752 1611
rect 6786 1577 6808 1611
rect 6842 1577 6847 1611
rect 6747 1572 6847 1577
rect 7059 1611 7159 1619
rect 7059 1577 7064 1611
rect 7098 1577 7120 1611
rect 7154 1577 7159 1611
rect 7059 1572 7159 1577
rect 7395 1611 7551 1619
rect 7395 1577 7400 1611
rect 7434 1577 7456 1611
rect 7490 1577 7512 1611
rect 7546 1577 7551 1611
rect 7395 1572 7551 1577
rect 7899 1611 8111 1619
rect 7899 1577 7904 1611
rect 7938 1577 7960 1611
rect 7994 1577 8016 1611
rect 8050 1577 8072 1611
rect 8106 1577 8111 1611
rect 7899 1572 8111 1577
rect 8459 1611 8559 1619
rect 8459 1577 8464 1611
rect 8498 1577 8520 1611
rect 8554 1577 8559 1611
rect 8459 1572 8559 1577
rect 8771 1611 8871 1619
rect 8771 1577 8776 1611
rect 8810 1577 8832 1611
rect 8866 1577 8871 1611
rect 8771 1572 8871 1577
rect 9107 1611 9263 1619
rect 9107 1577 9112 1611
rect 9146 1577 9168 1611
rect 9202 1577 9224 1611
rect 9258 1577 9263 1611
rect 9107 1572 9263 1577
rect 9611 1611 9823 1619
rect 9611 1577 9616 1611
rect 9650 1577 9672 1611
rect 9706 1577 9728 1611
rect 9762 1577 9784 1611
rect 9818 1577 9823 1611
rect 9611 1572 9823 1577
rect 10171 1611 10271 1619
rect 10171 1577 10176 1611
rect 10210 1577 10232 1611
rect 10266 1577 10271 1611
rect 10171 1572 10271 1577
use cc_inv  cc_inv_5
timestamp 1637401559
transform -1 0 1712 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_4
timestamp 1637401559
transform -1 0 3424 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_2
timestamp 1637401559
transform -1 0 5136 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_3
timestamp 1637401559
transform -1 0 6848 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_1
timestamp 1637401559
transform -1 0 8560 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_0
timestamp 1637401559
transform -1 0 10272 0 -1 1619
box -76 -16 1748 1650
use cc_inv  cc_inv_10
timestamp 1637401559
transform 1 0 602 0 1 1819
box -76 -16 1748 1650
use cc_inv  cc_inv_9
timestamp 1637401559
transform 1 0 2314 0 1 1819
box -76 -16 1748 1650
use cc_inv  cc_inv_7
timestamp 1637401559
transform 1 0 4026 0 1 1819
box -76 -16 1748 1650
use cc_inv  cc_inv_8
timestamp 1637401559
transform 1 0 5738 0 1 1819
box -76 -16 1748 1650
use cc_inv  cc_inv_6
timestamp 1637401559
transform 1 0 7450 0 1 1819
box -76 -16 1748 1650
<< end >>
