magic
tech sky130A
timestamp 1637401633
<< pwell >>
rect 264 1834 876 1850
rect 9462 1834 10598 1850
rect 264 1666 10598 1834
<< psubdiff >>
rect 2309 3550 2320 3580
rect 2350 3550 2380 3580
rect 2410 3550 2440 3580
rect 2470 3550 2500 3580
rect 2530 3550 2541 3580
rect 5072 3550 5080 3580
rect 5110 3550 5118 3580
rect 5192 3550 5200 3580
rect 5230 3550 5238 3580
rect 5252 3550 5260 3580
rect 5290 3550 5298 3580
rect 7889 3550 7900 3580
rect 7930 3550 7960 3580
rect 7990 3550 8020 3580
rect 8050 3550 8080 3580
rect 8110 3550 8121 3580
rect 2299 -80 2310 -50
rect 2340 -80 2370 -50
rect 2400 -80 2430 -50
rect 2460 -80 2490 -50
rect 2520 -80 2531 -50
rect 5059 -80 5070 -50
rect 5100 -80 5130 -50
rect 5160 -80 5190 -50
rect 5220 -80 5250 -50
rect 5280 -80 5291 -50
rect 7879 -80 7890 -50
rect 7920 -80 7950 -50
rect 7980 -80 8010 -50
rect 8040 -80 8070 -50
rect 8100 -80 8111 -50
<< psubdiffcont >>
rect 2320 3550 2350 3580
rect 2380 3550 2410 3580
rect 2440 3550 2470 3580
rect 2500 3550 2530 3580
rect 5080 3550 5110 3580
rect 5200 3550 5230 3580
rect 5260 3550 5290 3580
rect 7900 3550 7930 3580
rect 7960 3550 7990 3580
rect 8020 3550 8050 3580
rect 8080 3550 8110 3580
rect 2310 -80 2340 -50
rect 2370 -80 2400 -50
rect 2430 -80 2460 -50
rect 2490 -80 2520 -50
rect 5070 -80 5100 -50
rect 5130 -80 5160 -50
rect 5190 -80 5220 -50
rect 5250 -80 5280 -50
rect 7890 -80 7920 -50
rect 7950 -80 7980 -50
rect 8010 -80 8040 -50
rect 8070 -80 8100 -50
<< locali >>
rect 2309 3550 2318 3580
rect 2352 3550 2378 3580
rect 2412 3550 2438 3580
rect 2472 3550 2498 3580
rect 2532 3550 2541 3580
rect 5072 3550 5078 3580
rect 5112 3550 5118 3580
rect 5192 3550 5198 3580
rect 5232 3550 5238 3580
rect 5252 3550 5258 3580
rect 5292 3550 5298 3580
rect 7889 3550 7898 3580
rect 7932 3550 7958 3580
rect 7992 3550 8018 3580
rect 8052 3550 8078 3580
rect 8112 3550 8121 3580
rect 2299 -80 2308 -50
rect 2342 -80 2368 -50
rect 2402 -80 2428 -50
rect 2462 -80 2488 -50
rect 2522 -80 2531 -50
rect 5059 -80 5068 -50
rect 5102 -80 5128 -50
rect 5162 -80 5188 -50
rect 5222 -80 5248 -50
rect 5282 -80 5291 -50
rect 7879 -80 7888 -50
rect 7922 -80 7948 -50
rect 7982 -80 8008 -50
rect 8042 -80 8068 -50
rect 8102 -80 8111 -50
<< viali >>
rect 2318 3580 2352 3582
rect 2378 3580 2412 3582
rect 2438 3580 2472 3582
rect 2498 3580 2532 3582
rect 5078 3580 5112 3582
rect 2318 3550 2320 3580
rect 2320 3550 2350 3580
rect 2350 3550 2352 3580
rect 2378 3550 2380 3580
rect 2380 3550 2410 3580
rect 2410 3550 2412 3580
rect 2438 3550 2440 3580
rect 2440 3550 2470 3580
rect 2470 3550 2472 3580
rect 2498 3550 2500 3580
rect 2500 3550 2530 3580
rect 2530 3550 2532 3580
rect 5078 3550 5080 3580
rect 5080 3550 5110 3580
rect 5110 3550 5112 3580
rect 2318 3548 2352 3550
rect 2378 3548 2412 3550
rect 2438 3548 2472 3550
rect 2498 3548 2532 3550
rect 5078 3548 5112 3550
rect 5138 3548 5172 3582
rect 5198 3580 5232 3582
rect 5258 3580 5292 3582
rect 7898 3580 7932 3582
rect 7958 3580 7992 3582
rect 8018 3580 8052 3582
rect 8078 3580 8112 3582
rect 5198 3550 5200 3580
rect 5200 3550 5230 3580
rect 5230 3550 5232 3580
rect 5258 3550 5260 3580
rect 5260 3550 5290 3580
rect 5290 3550 5292 3580
rect 7898 3550 7900 3580
rect 7900 3550 7930 3580
rect 7930 3550 7932 3580
rect 7958 3550 7960 3580
rect 7960 3550 7990 3580
rect 7990 3550 7992 3580
rect 8018 3550 8020 3580
rect 8020 3550 8050 3580
rect 8050 3550 8052 3580
rect 8078 3550 8080 3580
rect 8080 3550 8110 3580
rect 8110 3550 8112 3580
rect 5198 3548 5232 3550
rect 5258 3548 5292 3550
rect 7898 3548 7932 3550
rect 7958 3548 7992 3550
rect 8018 3548 8052 3550
rect 8078 3548 8112 3550
rect 2308 -50 2342 -48
rect 2368 -50 2402 -48
rect 2428 -50 2462 -48
rect 2488 -50 2522 -48
rect 5068 -50 5102 -48
rect 5128 -50 5162 -48
rect 5188 -50 5222 -48
rect 5248 -50 5282 -48
rect 7888 -50 7922 -48
rect 7948 -50 7982 -48
rect 8008 -50 8042 -48
rect 8068 -50 8102 -48
rect 2308 -80 2310 -50
rect 2310 -80 2340 -50
rect 2340 -80 2342 -50
rect 2368 -80 2370 -50
rect 2370 -80 2400 -50
rect 2400 -80 2402 -50
rect 2428 -80 2430 -50
rect 2430 -80 2460 -50
rect 2460 -80 2462 -50
rect 2488 -80 2490 -50
rect 2490 -80 2520 -50
rect 2520 -80 2522 -50
rect 5068 -80 5070 -50
rect 5070 -80 5100 -50
rect 5100 -80 5102 -50
rect 5128 -80 5130 -50
rect 5130 -80 5160 -50
rect 5160 -80 5162 -50
rect 5188 -80 5190 -50
rect 5190 -80 5220 -50
rect 5220 -80 5222 -50
rect 5248 -80 5250 -50
rect 5250 -80 5280 -50
rect 5280 -80 5282 -50
rect 7888 -80 7890 -50
rect 7890 -80 7920 -50
rect 7920 -80 7922 -50
rect 7948 -80 7950 -50
rect 7950 -80 7980 -50
rect 7980 -80 7982 -50
rect 8008 -80 8010 -50
rect 8010 -80 8040 -50
rect 8040 -80 8042 -50
rect 8068 -80 8070 -50
rect 8070 -80 8100 -50
rect 8100 -80 8102 -50
rect 2308 -82 2342 -80
rect 2368 -82 2402 -80
rect 2428 -82 2462 -80
rect 2488 -82 2522 -80
rect 5068 -82 5102 -80
rect 5128 -82 5162 -80
rect 5188 -82 5222 -80
rect 5248 -82 5282 -80
rect 7888 -82 7922 -80
rect 7948 -82 7982 -80
rect 8008 -82 8042 -80
rect 8068 -82 8102 -80
<< metal1 >>
rect 2309 3584 2541 3590
rect 2309 3546 2316 3584
rect 2354 3546 2376 3584
rect 2414 3546 2436 3584
rect 2474 3546 2496 3584
rect 2534 3546 2541 3584
rect 2309 3540 2541 3546
rect 5069 3584 5301 3590
rect 5069 3546 5076 3584
rect 5114 3546 5136 3584
rect 5174 3546 5196 3584
rect 5234 3546 5256 3584
rect 5294 3546 5301 3584
rect 5069 3540 5301 3546
rect 7889 3584 8121 3590
rect 7889 3546 7896 3584
rect 7934 3546 7956 3584
rect 7994 3546 8016 3584
rect 8054 3546 8076 3584
rect 8114 3546 8121 3584
rect 7889 3540 8121 3546
rect 9457 3462 9500 3469
rect 3711 3459 3749 3462
rect 3711 3427 3714 3459
rect 3746 3427 3749 3459
rect 3711 3424 3749 3427
rect 3783 3459 3821 3462
rect 3783 3427 3786 3459
rect 3818 3427 3821 3459
rect 3783 3424 3821 3427
rect 3855 3459 3893 3462
rect 3855 3427 3858 3459
rect 3890 3427 3893 3459
rect 3855 3424 3893 3427
rect 6473 3459 6511 3462
rect 6473 3427 6476 3459
rect 6508 3427 6511 3459
rect 6473 3424 6511 3427
rect 6545 3459 6583 3462
rect 6545 3427 6548 3459
rect 6580 3427 6583 3459
rect 6545 3424 6583 3427
rect 6625 3459 6663 3462
rect 6625 3427 6628 3459
rect 6660 3427 6663 3459
rect 6625 3424 6663 3427
rect 9279 3459 9317 3462
rect 9279 3427 9282 3459
rect 9314 3427 9317 3459
rect 9279 3424 9317 3427
rect 9351 3459 9389 3462
rect 9351 3427 9354 3459
rect 9386 3427 9389 3459
rect 9351 3424 9389 3427
rect 9421 3459 9500 3462
rect 9421 3427 9424 3459
rect 9456 3427 9500 3459
rect 9421 3424 9500 3427
rect 9457 3419 9500 3424
rect 1959 2284 2037 2334
rect 3671 2284 3749 2334
rect 5383 2284 5461 2334
rect 7095 2284 7173 2334
rect 8807 2284 8885 2334
rect 877 1166 955 1216
rect 2589 1166 2667 1216
rect 4301 1166 4379 1216
rect 6013 1166 6091 1216
rect 7725 1166 7803 1216
rect 9437 1166 9515 1216
rect 3726 73 3764 76
rect 3726 41 3729 73
rect 3761 41 3764 73
rect 3726 38 3764 41
rect 3797 73 3835 76
rect 3797 41 3800 73
rect 3832 41 3835 73
rect 3797 38 3835 41
rect 3869 73 3907 76
rect 3869 41 3872 73
rect 3904 41 3907 73
rect 3869 38 3907 41
rect 6523 73 6561 76
rect 6523 41 6526 73
rect 6558 41 6561 73
rect 6523 38 6561 41
rect 6603 73 6641 76
rect 6603 41 6606 73
rect 6638 41 6641 73
rect 6603 38 6641 41
rect 6675 73 6713 76
rect 6675 41 6678 73
rect 6710 41 6713 73
rect 6675 38 6713 41
rect 9293 73 9331 76
rect 9293 41 9296 73
rect 9328 41 9331 73
rect 9293 38 9331 41
rect 9365 73 9403 76
rect 9365 41 9368 73
rect 9400 41 9403 73
rect 9365 38 9403 41
rect 9437 73 9475 76
rect 9437 41 9440 73
rect 9472 41 9475 73
rect 9437 38 9475 41
rect 2299 -46 2531 -40
rect 2299 -84 2306 -46
rect 2344 -84 2366 -46
rect 2404 -84 2426 -46
rect 2464 -84 2486 -46
rect 2524 -84 2531 -46
rect 2299 -90 2531 -84
rect 5059 -46 5291 -40
rect 5059 -84 5066 -46
rect 5104 -84 5126 -46
rect 5164 -84 5186 -46
rect 5224 -84 5246 -46
rect 5284 -84 5291 -46
rect 5059 -90 5291 -84
rect 7879 -46 8111 -40
rect 7879 -84 7886 -46
rect 7924 -84 7946 -46
rect 7984 -84 8006 -46
rect 8044 -84 8066 -46
rect 8104 -84 8111 -46
rect 7879 -90 8111 -84
<< via1 >>
rect 2316 3582 2354 3584
rect 2316 3548 2318 3582
rect 2318 3548 2352 3582
rect 2352 3548 2354 3582
rect 2316 3546 2354 3548
rect 2376 3582 2414 3584
rect 2376 3548 2378 3582
rect 2378 3548 2412 3582
rect 2412 3548 2414 3582
rect 2376 3546 2414 3548
rect 2436 3582 2474 3584
rect 2436 3548 2438 3582
rect 2438 3548 2472 3582
rect 2472 3548 2474 3582
rect 2436 3546 2474 3548
rect 2496 3582 2534 3584
rect 2496 3548 2498 3582
rect 2498 3548 2532 3582
rect 2532 3548 2534 3582
rect 2496 3546 2534 3548
rect 5076 3582 5114 3584
rect 5076 3548 5078 3582
rect 5078 3548 5112 3582
rect 5112 3548 5114 3582
rect 5076 3546 5114 3548
rect 5136 3582 5174 3584
rect 5136 3548 5138 3582
rect 5138 3548 5172 3582
rect 5172 3548 5174 3582
rect 5136 3546 5174 3548
rect 5196 3582 5234 3584
rect 5196 3548 5198 3582
rect 5198 3548 5232 3582
rect 5232 3548 5234 3582
rect 5196 3546 5234 3548
rect 5256 3582 5294 3584
rect 5256 3548 5258 3582
rect 5258 3548 5292 3582
rect 5292 3548 5294 3582
rect 5256 3546 5294 3548
rect 7896 3582 7934 3584
rect 7896 3548 7898 3582
rect 7898 3548 7932 3582
rect 7932 3548 7934 3582
rect 7896 3546 7934 3548
rect 7956 3582 7994 3584
rect 7956 3548 7958 3582
rect 7958 3548 7992 3582
rect 7992 3548 7994 3582
rect 7956 3546 7994 3548
rect 8016 3582 8054 3584
rect 8016 3548 8018 3582
rect 8018 3548 8052 3582
rect 8052 3548 8054 3582
rect 8016 3546 8054 3548
rect 8076 3582 8114 3584
rect 8076 3548 8078 3582
rect 8078 3548 8112 3582
rect 8112 3548 8114 3582
rect 8076 3546 8114 3548
rect 909 3427 941 3459
rect 980 3427 1012 3459
rect 1052 3427 1084 3459
rect 3714 3427 3746 3459
rect 3786 3427 3818 3459
rect 3858 3427 3890 3459
rect 6476 3427 6508 3459
rect 6548 3427 6580 3459
rect 6628 3427 6660 3459
rect 9282 3427 9314 3459
rect 9354 3427 9386 3459
rect 9424 3427 9456 3459
rect 880 41 912 73
rect 958 41 990 73
rect 1030 41 1062 73
rect 3729 41 3761 73
rect 3800 41 3832 73
rect 3872 41 3904 73
rect 6526 41 6558 73
rect 6606 41 6638 73
rect 6678 41 6710 73
rect 9296 41 9328 73
rect 9368 41 9400 73
rect 9440 41 9472 73
rect 2306 -48 2344 -46
rect 2306 -82 2308 -48
rect 2308 -82 2342 -48
rect 2342 -82 2344 -48
rect 2306 -84 2344 -82
rect 2366 -48 2404 -46
rect 2366 -82 2368 -48
rect 2368 -82 2402 -48
rect 2402 -82 2404 -48
rect 2366 -84 2404 -82
rect 2426 -48 2464 -46
rect 2426 -82 2428 -48
rect 2428 -82 2462 -48
rect 2462 -82 2464 -48
rect 2426 -84 2464 -82
rect 2486 -48 2524 -46
rect 2486 -82 2488 -48
rect 2488 -82 2522 -48
rect 2522 -82 2524 -48
rect 2486 -84 2524 -82
rect 5066 -48 5104 -46
rect 5066 -82 5068 -48
rect 5068 -82 5102 -48
rect 5102 -82 5104 -48
rect 5066 -84 5104 -82
rect 5126 -48 5164 -46
rect 5126 -82 5128 -48
rect 5128 -82 5162 -48
rect 5162 -82 5164 -48
rect 5126 -84 5164 -82
rect 5186 -48 5224 -46
rect 5186 -82 5188 -48
rect 5188 -82 5222 -48
rect 5222 -82 5224 -48
rect 5186 -84 5224 -82
rect 5246 -48 5284 -46
rect 5246 -82 5248 -48
rect 5248 -82 5282 -48
rect 5282 -82 5284 -48
rect 5246 -84 5284 -82
rect 7886 -48 7924 -46
rect 7886 -82 7888 -48
rect 7888 -82 7922 -48
rect 7922 -82 7924 -48
rect 7886 -84 7924 -82
rect 7946 -48 7984 -46
rect 7946 -82 7948 -48
rect 7948 -82 7982 -48
rect 7982 -82 7984 -48
rect 7946 -84 7984 -82
rect 8006 -48 8044 -46
rect 8006 -82 8008 -48
rect 8008 -82 8042 -48
rect 8042 -82 8044 -48
rect 8006 -84 8044 -82
rect 8066 -48 8104 -46
rect 8066 -82 8068 -48
rect 8068 -82 8102 -48
rect 8102 -82 8104 -48
rect 8066 -84 8104 -82
<< metal2 >>
rect 2309 3586 2541 3590
rect 2309 3544 2314 3586
rect 2356 3544 2374 3586
rect 2416 3544 2434 3586
rect 2476 3544 2494 3586
rect 2536 3544 2541 3586
rect 2309 3540 2541 3544
rect 5069 3586 5301 3590
rect 5069 3544 5074 3586
rect 5116 3544 5134 3586
rect 5176 3544 5194 3586
rect 5236 3544 5254 3586
rect 5296 3544 5301 3586
rect 5069 3540 5301 3544
rect 7889 3586 8121 3590
rect 7889 3544 7894 3586
rect 7936 3544 7954 3586
rect 7996 3544 8014 3586
rect 8056 3544 8074 3586
rect 8116 3544 8121 3586
rect 7889 3540 8121 3544
rect 902 3461 948 3466
rect 902 3425 907 3461
rect 943 3425 948 3461
rect 902 3420 948 3425
rect 973 3461 1019 3466
rect 973 3425 978 3461
rect 1014 3425 1019 3461
rect 973 3420 1019 3425
rect 1045 3461 1091 3466
rect 1045 3425 1050 3461
rect 1086 3425 1091 3461
rect 1045 3420 1091 3425
rect 3707 3461 3753 3466
rect 3707 3425 3712 3461
rect 3748 3425 3753 3461
rect 3707 3420 3753 3425
rect 3779 3461 3825 3466
rect 3779 3425 3784 3461
rect 3820 3425 3825 3461
rect 3779 3420 3825 3425
rect 3851 3461 3897 3466
rect 3851 3425 3856 3461
rect 3892 3425 3897 3461
rect 3851 3420 3897 3425
rect 6469 3461 6515 3466
rect 6469 3425 6474 3461
rect 6510 3425 6515 3461
rect 6469 3420 6515 3425
rect 6541 3461 6587 3466
rect 6541 3425 6546 3461
rect 6582 3425 6587 3461
rect 6541 3420 6587 3425
rect 6621 3461 6667 3466
rect 6621 3425 6626 3461
rect 6662 3425 6667 3461
rect 6621 3420 6667 3425
rect 9275 3461 9321 3466
rect 9275 3425 9280 3461
rect 9316 3425 9321 3461
rect 9275 3420 9321 3425
rect 9347 3461 9393 3466
rect 9347 3425 9352 3461
rect 9388 3425 9393 3461
rect 9347 3420 9393 3425
rect 9417 3461 9463 3466
rect 9417 3425 9422 3461
rect 9458 3425 9463 3461
rect 9417 3420 9463 3425
rect 873 75 919 80
rect 873 39 878 75
rect 914 39 919 75
rect 873 34 919 39
rect 951 75 997 80
rect 951 39 956 75
rect 992 39 997 75
rect 951 34 997 39
rect 1023 75 1069 80
rect 1023 39 1028 75
rect 1064 39 1069 75
rect 1023 34 1069 39
rect 3722 75 3768 80
rect 3722 39 3727 75
rect 3763 39 3768 75
rect 3722 34 3768 39
rect 3793 75 3839 80
rect 3793 39 3798 75
rect 3834 39 3839 75
rect 3793 34 3839 39
rect 3865 75 3911 80
rect 3865 39 3870 75
rect 3906 39 3911 75
rect 3865 34 3911 39
rect 6519 75 6565 80
rect 6519 39 6524 75
rect 6560 39 6565 75
rect 6519 34 6565 39
rect 6599 75 6645 80
rect 6599 39 6604 75
rect 6640 39 6645 75
rect 6599 34 6645 39
rect 6671 75 6717 80
rect 6671 39 6676 75
rect 6712 39 6717 75
rect 6671 34 6717 39
rect 9289 75 9335 80
rect 9289 39 9294 75
rect 9330 39 9335 75
rect 9289 34 9335 39
rect 9361 75 9407 80
rect 9361 39 9366 75
rect 9402 39 9407 75
rect 9361 34 9407 39
rect 9433 75 9479 80
rect 9433 39 9438 75
rect 9474 39 9479 75
rect 9433 34 9479 39
rect 2299 -44 2531 -40
rect 2299 -86 2304 -44
rect 2346 -86 2364 -44
rect 2406 -86 2424 -44
rect 2466 -86 2484 -44
rect 2526 -86 2531 -44
rect 2299 -90 2531 -86
rect 5059 -44 5291 -40
rect 5059 -86 5064 -44
rect 5106 -86 5124 -44
rect 5166 -86 5184 -44
rect 5226 -86 5244 -44
rect 5286 -86 5291 -44
rect 5059 -90 5291 -86
rect 7879 -44 8111 -40
rect 7879 -86 7884 -44
rect 7926 -86 7944 -44
rect 7986 -86 8004 -44
rect 8046 -86 8064 -44
rect 8106 -86 8111 -44
rect 7879 -90 8111 -86
<< via2 >>
rect 2314 3584 2356 3586
rect 2314 3546 2316 3584
rect 2316 3546 2354 3584
rect 2354 3546 2356 3584
rect 2314 3544 2356 3546
rect 2374 3584 2416 3586
rect 2374 3546 2376 3584
rect 2376 3546 2414 3584
rect 2414 3546 2416 3584
rect 2374 3544 2416 3546
rect 2434 3584 2476 3586
rect 2434 3546 2436 3584
rect 2436 3546 2474 3584
rect 2474 3546 2476 3584
rect 2434 3544 2476 3546
rect 2494 3584 2536 3586
rect 2494 3546 2496 3584
rect 2496 3546 2534 3584
rect 2534 3546 2536 3584
rect 2494 3544 2536 3546
rect 5074 3584 5116 3586
rect 5074 3546 5076 3584
rect 5076 3546 5114 3584
rect 5114 3546 5116 3584
rect 5074 3544 5116 3546
rect 5134 3584 5176 3586
rect 5134 3546 5136 3584
rect 5136 3546 5174 3584
rect 5174 3546 5176 3584
rect 5134 3544 5176 3546
rect 5194 3584 5236 3586
rect 5194 3546 5196 3584
rect 5196 3546 5234 3584
rect 5234 3546 5236 3584
rect 5194 3544 5236 3546
rect 5254 3584 5296 3586
rect 5254 3546 5256 3584
rect 5256 3546 5294 3584
rect 5294 3546 5296 3584
rect 5254 3544 5296 3546
rect 7894 3584 7936 3586
rect 7894 3546 7896 3584
rect 7896 3546 7934 3584
rect 7934 3546 7936 3584
rect 7894 3544 7936 3546
rect 7954 3584 7996 3586
rect 7954 3546 7956 3584
rect 7956 3546 7994 3584
rect 7994 3546 7996 3584
rect 7954 3544 7996 3546
rect 8014 3584 8056 3586
rect 8014 3546 8016 3584
rect 8016 3546 8054 3584
rect 8054 3546 8056 3584
rect 8014 3544 8056 3546
rect 8074 3584 8116 3586
rect 8074 3546 8076 3584
rect 8076 3546 8114 3584
rect 8114 3546 8116 3584
rect 8074 3544 8116 3546
rect 907 3459 943 3461
rect 907 3427 909 3459
rect 909 3427 941 3459
rect 941 3427 943 3459
rect 907 3425 943 3427
rect 978 3459 1014 3461
rect 978 3427 980 3459
rect 980 3427 1012 3459
rect 1012 3427 1014 3459
rect 978 3425 1014 3427
rect 1050 3459 1086 3461
rect 1050 3427 1052 3459
rect 1052 3427 1084 3459
rect 1084 3427 1086 3459
rect 1050 3425 1086 3427
rect 3712 3459 3748 3461
rect 3712 3427 3714 3459
rect 3714 3427 3746 3459
rect 3746 3427 3748 3459
rect 3712 3425 3748 3427
rect 3784 3459 3820 3461
rect 3784 3427 3786 3459
rect 3786 3427 3818 3459
rect 3818 3427 3820 3459
rect 3784 3425 3820 3427
rect 3856 3459 3892 3461
rect 3856 3427 3858 3459
rect 3858 3427 3890 3459
rect 3890 3427 3892 3459
rect 3856 3425 3892 3427
rect 6474 3459 6510 3461
rect 6474 3427 6476 3459
rect 6476 3427 6508 3459
rect 6508 3427 6510 3459
rect 6474 3425 6510 3427
rect 6546 3459 6582 3461
rect 6546 3427 6548 3459
rect 6548 3427 6580 3459
rect 6580 3427 6582 3459
rect 6546 3425 6582 3427
rect 6626 3459 6662 3461
rect 6626 3427 6628 3459
rect 6628 3427 6660 3459
rect 6660 3427 6662 3459
rect 6626 3425 6662 3427
rect 9280 3459 9316 3461
rect 9280 3427 9282 3459
rect 9282 3427 9314 3459
rect 9314 3427 9316 3459
rect 9280 3425 9316 3427
rect 9352 3459 9388 3461
rect 9352 3427 9354 3459
rect 9354 3427 9386 3459
rect 9386 3427 9388 3459
rect 9352 3425 9388 3427
rect 9422 3459 9458 3461
rect 9422 3427 9424 3459
rect 9424 3427 9456 3459
rect 9456 3427 9458 3459
rect 9422 3425 9458 3427
rect 878 73 914 75
rect 878 41 880 73
rect 880 41 912 73
rect 912 41 914 73
rect 878 39 914 41
rect 956 73 992 75
rect 956 41 958 73
rect 958 41 990 73
rect 990 41 992 73
rect 956 39 992 41
rect 1028 73 1064 75
rect 1028 41 1030 73
rect 1030 41 1062 73
rect 1062 41 1064 73
rect 1028 39 1064 41
rect 3727 73 3763 75
rect 3727 41 3729 73
rect 3729 41 3761 73
rect 3761 41 3763 73
rect 3727 39 3763 41
rect 3798 73 3834 75
rect 3798 41 3800 73
rect 3800 41 3832 73
rect 3832 41 3834 73
rect 3798 39 3834 41
rect 3870 73 3906 75
rect 3870 41 3872 73
rect 3872 41 3904 73
rect 3904 41 3906 73
rect 3870 39 3906 41
rect 6524 73 6560 75
rect 6524 41 6526 73
rect 6526 41 6558 73
rect 6558 41 6560 73
rect 6524 39 6560 41
rect 6604 73 6640 75
rect 6604 41 6606 73
rect 6606 41 6638 73
rect 6638 41 6640 73
rect 6604 39 6640 41
rect 6676 73 6712 75
rect 6676 41 6678 73
rect 6678 41 6710 73
rect 6710 41 6712 73
rect 6676 39 6712 41
rect 9294 73 9330 75
rect 9294 41 9296 73
rect 9296 41 9328 73
rect 9328 41 9330 73
rect 9294 39 9330 41
rect 9366 73 9402 75
rect 9366 41 9368 73
rect 9368 41 9400 73
rect 9400 41 9402 73
rect 9366 39 9402 41
rect 9438 73 9474 75
rect 9438 41 9440 73
rect 9440 41 9472 73
rect 9472 41 9474 73
rect 9438 39 9474 41
rect 2304 -46 2346 -44
rect 2304 -84 2306 -46
rect 2306 -84 2344 -46
rect 2344 -84 2346 -46
rect 2304 -86 2346 -84
rect 2364 -46 2406 -44
rect 2364 -84 2366 -46
rect 2366 -84 2404 -46
rect 2404 -84 2406 -46
rect 2364 -86 2406 -84
rect 2424 -46 2466 -44
rect 2424 -84 2426 -46
rect 2426 -84 2464 -46
rect 2464 -84 2466 -46
rect 2424 -86 2466 -84
rect 2484 -46 2526 -44
rect 2484 -84 2486 -46
rect 2486 -84 2524 -46
rect 2524 -84 2526 -46
rect 2484 -86 2526 -84
rect 5064 -46 5106 -44
rect 5064 -84 5066 -46
rect 5066 -84 5104 -46
rect 5104 -84 5106 -46
rect 5064 -86 5106 -84
rect 5124 -46 5166 -44
rect 5124 -84 5126 -46
rect 5126 -84 5164 -46
rect 5164 -84 5166 -46
rect 5124 -86 5166 -84
rect 5184 -46 5226 -44
rect 5184 -84 5186 -46
rect 5186 -84 5224 -46
rect 5224 -84 5226 -46
rect 5184 -86 5226 -84
rect 5244 -46 5286 -44
rect 5244 -84 5246 -46
rect 5246 -84 5284 -46
rect 5284 -84 5286 -46
rect 5244 -86 5286 -84
rect 7884 -46 7926 -44
rect 7884 -84 7886 -46
rect 7886 -84 7924 -46
rect 7924 -84 7926 -46
rect 7884 -86 7926 -84
rect 7944 -46 7986 -44
rect 7944 -84 7946 -46
rect 7946 -84 7984 -46
rect 7984 -84 7986 -46
rect 7944 -86 7986 -84
rect 8004 -46 8046 -44
rect 8004 -84 8006 -46
rect 8006 -84 8044 -46
rect 8044 -84 8046 -46
rect 8004 -86 8046 -84
rect 8064 -46 8106 -44
rect 8064 -84 8066 -46
rect 8066 -84 8104 -46
rect 8104 -84 8106 -46
rect 8064 -86 8106 -84
<< metal3 >>
rect 2309 3588 2541 3590
rect 2309 3542 2312 3588
rect 2358 3542 2372 3588
rect 2418 3542 2432 3588
rect 2478 3542 2492 3588
rect 2538 3542 2541 3588
rect 2309 3540 2541 3542
rect 5069 3588 5301 3590
rect 5069 3542 5072 3588
rect 5118 3542 5132 3588
rect 5178 3542 5192 3588
rect 5238 3542 5252 3588
rect 5298 3542 5301 3588
rect 5069 3540 5301 3542
rect 7889 3588 8121 3590
rect 7889 3542 7892 3588
rect 7938 3542 7952 3588
rect 7998 3542 8012 3588
rect 8058 3542 8072 3588
rect 8118 3542 8121 3588
rect 7889 3540 8121 3542
rect 900 3466 1085 3469
rect 900 3463 1091 3466
rect 900 3423 905 3463
rect 945 3423 976 3463
rect 1016 3423 1048 3463
rect 1088 3423 1091 3463
rect 900 3420 1091 3423
rect 3706 3463 3898 3469
rect 3706 3423 3710 3463
rect 3750 3423 3782 3463
rect 3822 3423 3854 3463
rect 3894 3423 3898 3463
rect 900 3419 1085 3420
rect 3706 3419 3898 3423
rect 6468 3463 6668 3469
rect 6468 3423 6472 3463
rect 6512 3423 6544 3463
rect 6584 3423 6624 3463
rect 6664 3423 6668 3463
rect 6468 3419 6668 3423
rect 9274 3463 9466 3469
rect 9274 3423 9278 3463
rect 9318 3423 9350 3463
rect 9390 3423 9420 3463
rect 9460 3423 9466 3463
rect 9274 3419 9466 3423
rect 873 77 1069 81
rect 873 37 876 77
rect 916 37 954 77
rect 994 37 1026 77
rect 1066 37 1069 77
rect 873 31 1069 37
rect 3721 77 3913 81
rect 3721 37 3725 77
rect 3765 37 3796 77
rect 3836 37 3868 77
rect 3908 37 3913 77
rect 3721 31 3913 37
rect 6518 77 6718 81
rect 6518 37 6522 77
rect 6562 37 6602 77
rect 6642 37 6674 77
rect 6714 37 6718 77
rect 6518 31 6718 37
rect 9288 77 9480 81
rect 9288 37 9292 77
rect 9332 37 9364 77
rect 9404 37 9436 77
rect 9476 37 9480 77
rect 9288 31 9480 37
rect 2299 -42 2531 -40
rect 2299 -88 2302 -42
rect 2348 -88 2362 -42
rect 2408 -88 2422 -42
rect 2468 -88 2482 -42
rect 2528 -88 2531 -42
rect 2299 -90 2531 -88
rect 5059 -42 5291 -40
rect 5059 -88 5062 -42
rect 5108 -88 5122 -42
rect 5168 -88 5182 -42
rect 5228 -88 5242 -42
rect 5288 -88 5291 -42
rect 5059 -90 5291 -88
rect 7879 -42 8111 -40
rect 7879 -88 7882 -42
rect 7928 -88 7942 -42
rect 7988 -88 8002 -42
rect 8048 -88 8062 -42
rect 8108 -88 8111 -42
rect 7879 -90 8111 -88
<< via3 >>
rect 2312 3586 2358 3588
rect 2312 3544 2314 3586
rect 2314 3544 2356 3586
rect 2356 3544 2358 3586
rect 2312 3542 2358 3544
rect 2372 3586 2418 3588
rect 2372 3544 2374 3586
rect 2374 3544 2416 3586
rect 2416 3544 2418 3586
rect 2372 3542 2418 3544
rect 2432 3586 2478 3588
rect 2432 3544 2434 3586
rect 2434 3544 2476 3586
rect 2476 3544 2478 3586
rect 2432 3542 2478 3544
rect 2492 3586 2538 3588
rect 2492 3544 2494 3586
rect 2494 3544 2536 3586
rect 2536 3544 2538 3586
rect 2492 3542 2538 3544
rect 5072 3586 5118 3588
rect 5072 3544 5074 3586
rect 5074 3544 5116 3586
rect 5116 3544 5118 3586
rect 5072 3542 5118 3544
rect 5132 3586 5178 3588
rect 5132 3544 5134 3586
rect 5134 3544 5176 3586
rect 5176 3544 5178 3586
rect 5132 3542 5178 3544
rect 5192 3586 5238 3588
rect 5192 3544 5194 3586
rect 5194 3544 5236 3586
rect 5236 3544 5238 3586
rect 5192 3542 5238 3544
rect 5252 3586 5298 3588
rect 5252 3544 5254 3586
rect 5254 3544 5296 3586
rect 5296 3544 5298 3586
rect 5252 3542 5298 3544
rect 7892 3586 7938 3588
rect 7892 3544 7894 3586
rect 7894 3544 7936 3586
rect 7936 3544 7938 3586
rect 7892 3542 7938 3544
rect 7952 3586 7998 3588
rect 7952 3544 7954 3586
rect 7954 3544 7996 3586
rect 7996 3544 7998 3586
rect 7952 3542 7998 3544
rect 8012 3586 8058 3588
rect 8012 3544 8014 3586
rect 8014 3544 8056 3586
rect 8056 3544 8058 3586
rect 8012 3542 8058 3544
rect 8072 3586 8118 3588
rect 8072 3544 8074 3586
rect 8074 3544 8116 3586
rect 8116 3544 8118 3586
rect 8072 3542 8118 3544
rect 905 3461 945 3463
rect 905 3425 907 3461
rect 907 3425 943 3461
rect 943 3425 945 3461
rect 905 3423 945 3425
rect 976 3461 1016 3463
rect 976 3425 978 3461
rect 978 3425 1014 3461
rect 1014 3425 1016 3461
rect 976 3423 1016 3425
rect 1048 3461 1088 3463
rect 1048 3425 1050 3461
rect 1050 3425 1086 3461
rect 1086 3425 1088 3461
rect 1048 3423 1088 3425
rect 3710 3461 3750 3463
rect 3710 3425 3712 3461
rect 3712 3425 3748 3461
rect 3748 3425 3750 3461
rect 3710 3423 3750 3425
rect 3782 3461 3822 3463
rect 3782 3425 3784 3461
rect 3784 3425 3820 3461
rect 3820 3425 3822 3461
rect 3782 3423 3822 3425
rect 3854 3461 3894 3463
rect 3854 3425 3856 3461
rect 3856 3425 3892 3461
rect 3892 3425 3894 3461
rect 3854 3423 3894 3425
rect 6472 3461 6512 3463
rect 6472 3425 6474 3461
rect 6474 3425 6510 3461
rect 6510 3425 6512 3461
rect 6472 3423 6512 3425
rect 6544 3461 6584 3463
rect 6544 3425 6546 3461
rect 6546 3425 6582 3461
rect 6582 3425 6584 3461
rect 6544 3423 6584 3425
rect 6624 3461 6664 3463
rect 6624 3425 6626 3461
rect 6626 3425 6662 3461
rect 6662 3425 6664 3461
rect 6624 3423 6664 3425
rect 9278 3461 9318 3463
rect 9278 3425 9280 3461
rect 9280 3425 9316 3461
rect 9316 3425 9318 3461
rect 9278 3423 9318 3425
rect 9350 3461 9390 3463
rect 9350 3425 9352 3461
rect 9352 3425 9388 3461
rect 9388 3425 9390 3461
rect 9350 3423 9390 3425
rect 9420 3461 9460 3463
rect 9420 3425 9422 3461
rect 9422 3425 9458 3461
rect 9458 3425 9460 3461
rect 9420 3423 9460 3425
rect 876 75 916 77
rect 876 39 878 75
rect 878 39 914 75
rect 914 39 916 75
rect 876 37 916 39
rect 954 75 994 77
rect 954 39 956 75
rect 956 39 992 75
rect 992 39 994 75
rect 954 37 994 39
rect 1026 75 1066 77
rect 1026 39 1028 75
rect 1028 39 1064 75
rect 1064 39 1066 75
rect 1026 37 1066 39
rect 3725 75 3765 77
rect 3725 39 3727 75
rect 3727 39 3763 75
rect 3763 39 3765 75
rect 3725 37 3765 39
rect 3796 75 3836 77
rect 3796 39 3798 75
rect 3798 39 3834 75
rect 3834 39 3836 75
rect 3796 37 3836 39
rect 3868 75 3908 77
rect 3868 39 3870 75
rect 3870 39 3906 75
rect 3906 39 3908 75
rect 3868 37 3908 39
rect 6522 75 6562 77
rect 6522 39 6524 75
rect 6524 39 6560 75
rect 6560 39 6562 75
rect 6522 37 6562 39
rect 6602 75 6642 77
rect 6602 39 6604 75
rect 6604 39 6640 75
rect 6640 39 6642 75
rect 6602 37 6642 39
rect 6674 75 6714 77
rect 6674 39 6676 75
rect 6676 39 6712 75
rect 6712 39 6714 75
rect 6674 37 6714 39
rect 9292 75 9332 77
rect 9292 39 9294 75
rect 9294 39 9330 75
rect 9330 39 9332 75
rect 9292 37 9332 39
rect 9364 75 9404 77
rect 9364 39 9366 75
rect 9366 39 9402 75
rect 9402 39 9404 75
rect 9364 37 9404 39
rect 9436 75 9476 77
rect 9436 39 9438 75
rect 9438 39 9474 75
rect 9474 39 9476 75
rect 9436 37 9476 39
rect 2302 -44 2348 -42
rect 2302 -86 2304 -44
rect 2304 -86 2346 -44
rect 2346 -86 2348 -44
rect 2302 -88 2348 -86
rect 2362 -44 2408 -42
rect 2362 -86 2364 -44
rect 2364 -86 2406 -44
rect 2406 -86 2408 -44
rect 2362 -88 2408 -86
rect 2422 -44 2468 -42
rect 2422 -86 2424 -44
rect 2424 -86 2466 -44
rect 2466 -86 2468 -44
rect 2422 -88 2468 -86
rect 2482 -44 2528 -42
rect 2482 -86 2484 -44
rect 2484 -86 2526 -44
rect 2526 -86 2528 -44
rect 2482 -88 2528 -86
rect 5062 -44 5108 -42
rect 5062 -86 5064 -44
rect 5064 -86 5106 -44
rect 5106 -86 5108 -44
rect 5062 -88 5108 -86
rect 5122 -44 5168 -42
rect 5122 -86 5124 -44
rect 5124 -86 5166 -44
rect 5166 -86 5168 -44
rect 5122 -88 5168 -86
rect 5182 -44 5228 -42
rect 5182 -86 5184 -44
rect 5184 -86 5226 -44
rect 5226 -86 5228 -44
rect 5182 -88 5228 -86
rect 5242 -44 5288 -42
rect 5242 -86 5244 -44
rect 5244 -86 5286 -44
rect 5286 -86 5288 -44
rect 5242 -88 5288 -86
rect 7882 -44 7928 -42
rect 7882 -86 7884 -44
rect 7884 -86 7926 -44
rect 7926 -86 7928 -44
rect 7882 -88 7928 -86
rect 7942 -44 7988 -42
rect 7942 -86 7944 -44
rect 7944 -86 7986 -44
rect 7986 -86 7988 -44
rect 7942 -88 7988 -86
rect 8002 -44 8048 -42
rect 8002 -86 8004 -44
rect 8004 -86 8046 -44
rect 8046 -86 8048 -44
rect 8002 -88 8048 -86
rect 8062 -44 8108 -42
rect 8062 -86 8064 -44
rect 8064 -86 8106 -44
rect 8106 -86 8108 -44
rect 8062 -88 8108 -86
<< metal4 >>
rect 2309 3588 2541 3590
rect 2309 3542 2312 3588
rect 2358 3542 2372 3588
rect 2418 3542 2432 3588
rect 2478 3542 2492 3588
rect 2538 3542 2541 3588
rect 2309 3540 2541 3542
rect 5069 3588 5125 3590
rect 5069 3542 5072 3588
rect 5118 3542 5125 3588
rect 5069 3540 5125 3542
rect 5300 3540 5301 3590
rect 7889 3588 8121 3590
rect 7889 3542 7892 3588
rect 7938 3542 7952 3588
rect 7998 3542 8012 3588
rect 8058 3542 8072 3588
rect 8118 3542 8121 3588
rect 7889 3540 8121 3542
rect 3706 3463 3754 3469
rect 3706 3423 3710 3463
rect 3750 3423 3754 3463
rect 3706 3419 3754 3423
rect 3778 3463 3826 3469
rect 3778 3423 3782 3463
rect 3822 3423 3826 3463
rect 3778 3419 3826 3423
rect 3850 3463 3898 3469
rect 3850 3423 3854 3463
rect 3894 3423 3898 3463
rect 3850 3419 3898 3423
rect 6468 3463 6516 3469
rect 6468 3423 6472 3463
rect 6512 3423 6516 3463
rect 6468 3419 6516 3423
rect 6540 3463 6588 3469
rect 6540 3423 6544 3463
rect 6584 3423 6588 3463
rect 6540 3419 6588 3423
rect 6620 3463 6668 3469
rect 6620 3423 6624 3463
rect 6664 3423 6668 3463
rect 6620 3419 6668 3423
rect 9274 3463 9322 3469
rect 9274 3423 9278 3463
rect 9318 3423 9322 3463
rect 9274 3419 9322 3423
rect 9346 3463 9394 3469
rect 9346 3423 9350 3463
rect 9390 3423 9394 3463
rect 9346 3419 9394 3423
rect 9416 3463 9464 3469
rect 9416 3423 9420 3463
rect 9460 3423 9464 3463
rect 9416 3419 9464 3423
rect 873 77 1069 81
rect 873 37 876 77
rect 916 37 954 77
rect 994 37 1026 77
rect 1066 37 1069 77
rect 873 31 1069 37
rect 3721 77 3769 81
rect 3721 37 3725 77
rect 3765 37 3769 77
rect 3721 31 3769 37
rect 3792 77 3840 81
rect 3792 37 3796 77
rect 3836 37 3840 77
rect 3792 31 3840 37
rect 3864 77 3912 81
rect 3864 37 3868 77
rect 3908 37 3912 77
rect 3864 31 3912 37
rect 6518 77 6566 81
rect 6518 37 6522 77
rect 6562 37 6566 77
rect 6518 31 6566 37
rect 6598 77 6646 81
rect 6598 37 6602 77
rect 6642 37 6646 77
rect 6598 31 6646 37
rect 6670 77 6718 81
rect 6670 37 6674 77
rect 6714 37 6718 77
rect 6670 31 6718 37
rect 9288 77 9336 81
rect 9288 37 9292 77
rect 9332 37 9336 77
rect 9288 31 9336 37
rect 9360 77 9408 81
rect 9360 37 9364 77
rect 9404 37 9408 77
rect 9360 31 9408 37
rect 9432 77 9480 81
rect 9432 37 9436 77
rect 9476 37 9480 77
rect 9432 31 9480 37
rect 2299 -42 2531 -40
rect 2299 -88 2302 -42
rect 2348 -88 2362 -42
rect 2408 -88 2422 -42
rect 2468 -88 2482 -42
rect 2528 -88 2531 -42
rect 2299 -90 2531 -88
rect 5059 -42 5291 -40
rect 5059 -88 5062 -42
rect 5108 -88 5122 -42
rect 5168 -88 5182 -42
rect 5228 -88 5242 -42
rect 5288 -88 5291 -42
rect 5059 -90 5291 -88
rect 7879 -42 8111 -40
rect 7879 -88 7882 -42
rect 7928 -88 7942 -42
rect 7988 -88 8002 -42
rect 8048 -88 8062 -42
rect 8108 -88 8111 -42
rect 7879 -90 8111 -88
use ring_osc  ring_osc_0
timestamp 1637401559
transform 1 0 300 0 1 31
box -300 -31 10550 3469
use pwell_co_ring  pwell_co_ring_0
timestamp 1637401559
transform 1 0 170 0 1 -80
box 0 0 10560 3660
use power_ring  power_ring_0
timestamp 1637401559
transform 1 0 -900 0 1 -3500
box 0 0 12200 10500
<< labels >>
flabel metal1 912 1191 912 1191 1 FreeSans 800 0 0 0 p[0]
port 1 s signal output
flabel metal1 2624 1191 2624 1191 1 FreeSans 800 0 0 0 p[2]
port 3 s signal output
flabel metal1 4336 1191 4336 1191 1 FreeSans 800 0 0 0 p[4]
port 5 s signal output
flabel metal1 6048 1191 6048 1191 1 FreeSans 800 0 0 0 p[6]
port 7 s signal output
flabel metal1 7760 1191 7760 1191 1 FreeSans 800 0 0 0 p[8]
port 9 s signal output
flabel metal1 9472 1191 9472 1191 1 FreeSans 800 0 0 0 p[10]
port 11 s signal output
flabel metal1 2002 2309 2002 2309 1 FreeSans 800 0 0 0 p[1]
port 2 s signal output
flabel metal1 3714 2309 3714 2309 1 FreeSans 800 0 0 0 p[3]
port 4 s signal output
flabel metal1 5426 2309 5426 2309 1 FreeSans 800 0 0 0 p[5]
port 6 s signal output
flabel metal1 7138 2309 7138 2309 1 FreeSans 800 0 0 0 p[7]
port 8 s signal output
flabel metal1 8850 2309 8850 2309 1 FreeSans 800 0 0 0 p[9]
port 10 s signal output
<< end >>
