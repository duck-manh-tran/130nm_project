magic
tech sky130A
timestamp 1623843753
<< locali >>
rect -540 2428 -500 2430
rect -540 2402 -538 2428
rect -512 2402 -500 2428
rect -540 2400 -500 2402
<< viali >>
rect -538 2402 -512 2428
<< obsli1 >>
rect -500 2480 11700 3100
rect -440 2350 11700 2480
rect -500 -120 11700 2350
<< metal1 >>
rect -545 2428 -505 2435
rect -545 2402 -538 2428
rect -512 2402 -505 2428
rect -545 2395 -505 2402
<< obsm1 >>
rect -500 2480 11700 3100
rect -440 2350 11700 2480
rect -500 -120 11700 2350
<< metal2 >>
rect 2208 3108 2250 3150
rect 4645 3108 4687 3150
rect 6324 3108 6366 3150
rect 7854 3108 7896 3150
rect 10097 3108 10139 3150
rect 11760 1900 11810 1950
rect 211 -172 253 -130
rect 2025 -172 2067 -130
rect 3800 -172 3842 -130
rect 6099 -172 6141 -130
rect 7431 -172 7473 -130
rect 9111 -172 9153 -130
<< obsm2 >>
rect -500 3050 2150 3100
rect 2310 3050 4580 3100
rect 4740 3050 6260 3100
rect 6420 3050 7796 3100
rect 7956 3050 9982 3100
rect -500 3012 9982 3050
rect 10235 3012 11752 3100
rect -500 2480 11752 3012
rect -440 2350 11752 2480
rect -500 2007 11752 2350
rect -500 1847 11702 2007
rect -500 -70 11752 1847
rect -500 -120 154 -70
rect 314 -120 1963 -70
rect 2123 -120 3740 -70
rect 3900 -120 6040 -70
rect 6200 -120 7371 -70
rect 7531 -120 9052 -70
rect 9212 -120 11752 -70
<< metal3 >>
rect -500 6500 2100 6700
rect 8800 -3400 11300 -3200
<< obsm3 >>
rect -500 2480 11700 3100
rect -440 2350 11700 2480
rect -500 -120 11700 2350
use power_ring  power_ring_0
timestamp 1623832439
transform 1 0 -500 0 1 -3800
box 0 0 12200 10500
<< labels >>
flabel metal1 -545 2395 -505 2435 1 FreeSans 8 0 0 0 enb
port 12 w signal input
flabel metal3 -500 6500 2100 6700 1 FreeSans 8 0 0 0 vccd2
port 14 n power bidirectional
flabel metal3 8800 -3400 11300 -3200 1 FreeSans 8 0 0 0 vssd2
port 15 s ground bidirectional
flabel metal2 2208 3108 2250 3150 1 FreeSans 8 0 0 0 p[6]
port 7 n signal output
flabel metal2 4645 3108 4687 3150 1 FreeSans 8 0 0 0 p[7]
port 8 n signal output
flabel metal2 6324 3108 6366 3150 1 FreeSans 8 0 0 0 p[8]
port 9 n signal output
flabel metal2 10097 3108 10139 3150 1 FreeSans 8 0 0 0 p[10]
port 11 n signal output
flabel metal2 9111 -172 9153 -130 1 FreeSans 8 0 0 0 p[0]
port 1 s signal output
flabel metal2 7431 -172 7473 -130 1 FreeSans 8 0 0 0 p[1]
port 2 s signal output
flabel metal2 6099 -172 6141 -130 1 FreeSans 8 0 0 0 p[2]
port 3 s signal output
flabel metal2 3800 -172 3842 -130 1 FreeSans 8 0 0 0 p[3]
port 4 s signal output
flabel metal2 2025 -172 2067 -130 1 FreeSans 8 0 0 0 p[4]
port 5 s signal output
flabel metal2 211 -172 253 -130 1 FreeSans 8 0 0 0 p[5]
port 6 s signal output
flabel metal2 7854 3108 7896 3150 1 FreeSans 8 0 0 0 p[9]
port 10 nsew default output
flabel metal2 11760 1900 11810 1950 1 FreeSans 8 0 0 0 input_analog
port 13 nsew signal input
<< end >>
