magic
tech sky130A
timestamp 1637149740
<< pwell >>
rect 209 598 226 610
rect 757 598 774 610
<< poly >>
rect 95 652 505 700
rect 95 635 101 652
rect 118 635 137 652
rect 154 635 173 652
rect 190 635 209 652
rect 226 635 374 652
rect 391 635 410 652
rect 427 635 446 652
rect 463 635 482 652
rect 499 635 505 652
rect 95 615 505 635
rect 95 598 101 615
rect 118 598 137 615
rect 154 598 173 615
rect 190 598 209 615
rect 226 598 374 615
rect 391 598 410 615
rect 427 598 446 615
rect 463 598 482 615
rect 499 598 505 615
rect 95 550 505 598
rect 643 652 1053 700
rect 643 635 649 652
rect 666 635 685 652
rect 702 635 721 652
rect 738 635 757 652
rect 774 635 922 652
rect 939 635 958 652
rect 975 635 994 652
rect 1011 635 1030 652
rect 1047 635 1053 652
rect 643 615 1053 635
rect 643 598 649 615
rect 666 598 685 615
rect 702 598 721 615
rect 738 598 757 615
rect 774 598 922 615
rect 939 598 958 615
rect 975 598 994 615
rect 1011 598 1030 615
rect 1047 598 1053 615
rect 643 550 1053 598
<< polycont >>
rect 101 635 118 652
rect 137 635 154 652
rect 173 635 190 652
rect 209 635 226 652
rect 374 635 391 652
rect 410 635 427 652
rect 446 635 463 652
rect 482 635 499 652
rect 101 598 118 615
rect 137 598 154 615
rect 173 598 190 615
rect 209 598 226 615
rect 374 598 391 615
rect 410 598 427 615
rect 446 598 463 615
rect 482 598 499 615
rect 649 635 666 652
rect 685 635 702 652
rect 721 635 738 652
rect 757 635 774 652
rect 922 635 939 652
rect 958 635 975 652
rect 994 635 1011 652
rect 1030 635 1047 652
rect 649 598 666 615
rect 685 598 702 615
rect 721 598 738 615
rect 757 598 774 615
rect 922 598 939 615
rect 958 598 975 615
rect 994 598 1011 615
rect 1030 598 1047 615
<< locali >>
rect 93 635 101 652
rect 118 635 137 652
rect 154 635 173 652
rect 190 635 209 652
rect 226 635 234 652
rect 93 598 101 615
rect 118 598 137 615
rect 154 598 173 615
rect 190 598 209 615
rect 226 598 234 615
rect 285 498 315 749
rect 366 635 374 652
rect 391 635 410 652
rect 427 635 446 652
rect 463 635 482 652
rect 499 635 507 652
rect 641 635 649 652
rect 666 635 685 652
rect 702 635 721 652
rect 738 635 757 652
rect 774 635 782 652
rect 366 598 374 615
rect 391 598 410 615
rect 427 598 446 615
rect 463 598 482 615
rect 499 598 507 615
rect 641 598 649 615
rect 666 598 685 615
rect 702 598 721 615
rect 738 598 757 615
rect 774 598 782 615
rect 833 498 863 749
rect 914 635 922 652
rect 939 635 958 652
rect 975 635 994 652
rect 1011 635 1030 652
rect 1047 635 1055 652
rect 914 598 922 615
rect 939 598 958 615
rect 975 598 994 615
rect 1011 598 1030 615
rect 1047 598 1055 615
rect 1845 451 1875 793
<< viali >>
rect 101 635 118 652
rect 137 635 154 652
rect 173 635 190 652
rect 209 635 226 652
rect 101 598 118 615
rect 137 598 154 615
rect 173 598 190 615
rect 209 598 226 615
rect 374 635 391 652
rect 410 635 427 652
rect 446 635 463 652
rect 482 635 499 652
rect 649 635 666 652
rect 685 635 702 652
rect 721 635 738 652
rect 757 635 774 652
rect 374 598 391 615
rect 410 598 427 615
rect 446 598 463 615
rect 482 598 499 615
rect 649 598 666 615
rect 685 598 702 615
rect 721 598 738 615
rect 757 598 774 615
rect 922 635 939 652
rect 958 635 975 652
rect 994 635 1011 652
rect 1030 635 1047 652
rect 922 598 939 615
rect 958 598 975 615
rect 994 598 1011 615
rect 1030 598 1047 615
<< metal1 >>
rect 95 652 234 655
rect 95 635 101 652
rect 118 635 137 652
rect 154 635 173 652
rect 190 635 209 652
rect 226 650 234 652
rect 366 652 505 655
rect 366 650 374 652
rect 226 635 374 650
rect 391 635 410 652
rect 427 635 446 652
rect 463 635 482 652
rect 499 635 505 652
rect 95 615 505 635
rect 95 598 101 615
rect 118 598 137 615
rect 154 598 173 615
rect 190 598 209 615
rect 226 600 374 615
rect 226 598 234 600
rect 95 595 234 598
rect 366 598 374 600
rect 391 598 410 615
rect 427 598 446 615
rect 463 598 482 615
rect 499 598 505 615
rect 366 595 505 598
rect 643 652 782 655
rect 643 635 649 652
rect 666 635 685 652
rect 702 635 721 652
rect 738 635 757 652
rect 774 650 782 652
rect 914 652 1053 655
rect 914 650 922 652
rect 774 635 922 650
rect 939 635 958 652
rect 975 635 994 652
rect 1011 635 1030 652
rect 1047 635 1053 652
rect 643 615 1053 635
rect 643 598 649 615
rect 666 598 685 615
rect 702 598 721 615
rect 738 598 757 615
rect 774 600 922 615
rect 774 598 782 600
rect 643 595 782 598
rect 914 598 922 600
rect 939 598 958 615
rect 975 598 994 615
rect 1011 598 1030 615
rect 1047 598 1053 615
rect 914 595 1053 598
use pfet_34  pfet_34_0
timestamp 1637141615
transform 1 0 1550 0 1 650
box 0 0 400 1000
use nfet_34  nfet_34_0
timestamp 1637142191
transform 1 0 1550 0 1 0
box 0 0 400 610
use pfet_12  pfet_12_1
timestamp 1637143825
transform 1 0 498 0 1 650
box 0 0 700 1000
use nfet_12  nfet_12_1
timestamp 1637148458
transform 1 0 548 0 1 0
box 0 0 600 610
use pfet_12  pfet_12_0
timestamp 1637143825
transform 1 0 -50 0 1 650
box 0 0 700 1000
use nfet_12  nfet_12_0
timestamp 1637148458
transform 1 0 0 0 1 0
box 0 0 600 610
<< end >>
