magic
tech sky130A
magscale 1 2
timestamp 1623122433
<< psubdiff >>
rect 3176 14400 3300 14500
rect 3400 14400 3500 14500
rect 3600 14400 3700 14500
rect 3800 14400 3900 14500
rect 4000 14400 4100 14500
rect 4200 14400 4300 14500
rect 4400 14400 4500 14500
rect 4600 14400 4700 14500
rect 4800 14400 4900 14500
rect 5000 14400 5100 14500
rect 5200 14400 5300 14500
rect 5400 14400 5500 14500
rect 5600 14400 5700 14500
rect 5800 14400 5900 14500
rect 6000 14400 6100 14500
rect 6200 14400 6300 14500
rect 6400 14400 6500 14500
rect 6600 14400 6700 14500
rect 6800 14400 6900 14500
rect 7000 14400 7100 14500
rect 7200 14400 7300 14500
rect 7400 14400 7500 14500
rect 7600 14400 7700 14500
rect 7800 14400 7900 14500
rect 8000 14400 8100 14500
rect 8200 14400 8300 14500
rect 8400 14400 8500 14500
rect 8600 14400 8700 14500
rect 8800 14400 8900 14500
rect 9000 14400 9100 14500
rect 9200 14400 9300 14500
rect 9400 14400 9500 14500
rect 9600 14400 9700 14500
rect 9800 14400 9900 14500
rect 10000 14400 10100 14500
rect 10200 14400 10300 14500
rect 10400 14400 10500 14500
rect 10600 14400 10700 14500
rect 10800 14400 10900 14500
rect 11000 14400 11100 14500
rect 11200 14400 11300 14500
rect 11400 14400 11500 14500
rect 11600 14400 11700 14500
rect 11800 14400 11900 14500
rect 12000 14400 12100 14500
rect 12200 14400 12300 14500
rect 12400 14400 12500 14500
rect 12600 14400 12700 14500
rect 12800 14400 12900 14500
rect 13000 14400 13100 14500
rect 13200 14400 13300 14500
rect 13400 14400 13500 14500
rect 13600 14400 13700 14500
rect 13800 14400 13900 14500
rect 14000 14400 14100 14500
rect 14200 14400 14300 14500
rect 14400 14400 14500 14500
rect 14600 14400 14700 14500
rect 14800 14400 14900 14500
rect 15000 14400 15100 14500
rect 15200 14400 15300 14500
rect 15400 14400 15500 14500
rect 15600 14400 15700 14500
rect 15800 14400 15900 14500
rect 16000 14400 16100 14500
rect 16200 14400 16300 14500
rect 16400 14400 16500 14500
rect 16600 14400 16700 14500
rect 16800 14400 16900 14500
rect 17000 14400 17100 14500
rect 17200 14400 17300 14500
rect 17400 14400 17500 14500
rect 17600 14400 17700 14500
rect 17800 14400 17900 14500
rect 18000 14400 18100 14500
rect 18200 14400 18300 14500
rect 18400 14400 18500 14500
rect 18600 14400 18700 14500
rect 18800 14400 18900 14500
rect 19000 14400 19100 14500
rect 19200 14400 19300 14500
rect 19400 14400 19500 14500
rect 19600 14400 19700 14500
rect 19800 14400 19900 14500
rect 20000 14400 20100 14500
rect 20200 14400 20300 14500
rect 20400 14400 20500 14500
rect 20600 14400 20700 14500
rect 20800 14400 20900 14500
rect 21000 14400 21100 14500
rect 21200 14400 21300 14500
rect 21400 14400 21500 14500
rect 21600 14400 21700 14500
rect 21800 14400 21900 14500
rect 22000 14400 22100 14500
rect 22200 14400 22300 14500
rect 22400 14400 22500 14500
rect 22600 14400 22700 14500
rect 22800 14400 22900 14500
rect 23000 14400 23100 14500
rect 23200 14400 23300 14500
rect 23400 14400 23500 14500
rect 23600 14400 23700 14500
rect 23800 14400 23900 14500
rect 24000 14400 24100 14500
rect 24200 14400 24300 14500
rect 24400 14400 24500 14500
rect 24600 14400 24700 14500
rect 24800 14400 24900 14500
rect 25000 14400 25100 14500
rect 25200 14400 25300 14500
rect 25400 14400 25500 14500
rect 25600 14400 25700 14500
rect 25800 14400 25900 14500
rect 26000 14400 26100 14500
rect 26200 14400 26300 14500
rect 26400 14400 26500 14500
rect 26600 14400 26700 14500
rect 26800 14400 26900 14500
rect 27000 14400 27100 14500
rect 27200 14400 27300 14500
rect 27400 14400 27500 14500
rect 27600 14400 27700 14500
rect 27800 14400 27900 14500
rect 28000 14400 28100 14500
rect 28200 14400 28300 14500
rect 28400 14400 28500 14500
rect 28600 14400 28700 14500
rect 28800 14400 28900 14500
rect 29000 14400 29100 14500
rect 29200 14400 29300 14500
rect 29400 14400 29500 14500
rect 29600 14400 29700 14500
rect 29800 14400 29900 14500
rect 30000 14400 30100 14500
rect 30200 14400 30300 14500
rect 30400 14400 30500 14500
rect 30600 14400 30700 14500
rect 30800 14400 30900 14500
rect 31000 14400 31100 14500
rect 31200 14400 31300 14500
rect 31400 14400 31500 14500
rect 31600 14400 31700 14500
rect 31800 14400 31900 14500
rect 32000 14400 32100 14500
rect 32200 14400 32300 14500
rect 32400 14400 32500 14500
rect 32600 14400 32700 14500
rect 32800 14400 32900 14500
rect 33000 14400 33100 14500
rect 33200 14400 33324 14500
rect 3200 14300 3300 14400
rect 3200 14100 3300 14200
rect 3200 13900 3300 14000
rect 3200 13700 3300 13800
rect 3200 13500 3300 13600
rect 3200 13300 3300 13400
rect 3200 13100 3300 13200
rect 3200 12900 3300 13000
rect 3200 12700 3300 12800
rect 3200 12500 3300 12600
rect 3200 12300 3300 12400
rect 3200 12100 3300 12200
rect 3200 11900 3300 12000
rect 3200 11700 3300 11800
rect 3200 11500 3300 11600
rect 3200 11300 3300 11400
rect 3200 11100 3300 11200
rect 3200 10900 3300 11000
rect 3200 10700 3300 10800
rect 3200 10500 3300 10600
rect 33200 14300 33300 14400
rect 33200 14100 33300 14200
rect 33200 13900 33300 14000
rect 33200 13700 33300 13800
rect 33200 13500 33300 13600
rect 33200 13300 33300 13400
rect 33200 13100 33300 13200
rect 33200 12900 33300 13000
rect 33200 12700 33300 12800
rect 33200 12500 33300 12600
rect 33200 12300 33300 12400
rect 33200 12100 33300 12200
rect 33200 11900 33300 12000
rect 33200 11700 33300 11800
rect 33200 11500 33300 11600
rect 33200 11300 33300 11400
rect 33200 11100 33300 11200
rect 33200 10900 33300 11000
rect 33200 10700 33300 10800
rect 33200 10500 33300 10600
rect 3176 10400 3300 10500
rect 3400 10400 3500 10500
rect 3600 10400 3700 10500
rect 3800 10400 3900 10500
rect 4000 10400 4100 10500
rect 4200 10400 4300 10500
rect 4400 10400 4500 10500
rect 4600 10400 4700 10500
rect 4800 10400 4900 10500
rect 5000 10400 5100 10500
rect 5200 10400 5300 10500
rect 5400 10400 5500 10500
rect 5600 10400 5700 10500
rect 5800 10400 5900 10500
rect 6000 10400 6100 10500
rect 6200 10400 6300 10500
rect 6400 10400 6500 10500
rect 6600 10400 6700 10500
rect 6800 10400 6900 10500
rect 7000 10400 7100 10500
rect 7200 10400 7300 10500
rect 7400 10400 7500 10500
rect 7600 10400 7700 10500
rect 7800 10400 7900 10500
rect 8000 10400 8100 10500
rect 8200 10400 8300 10500
rect 8400 10400 8500 10500
rect 8600 10400 8700 10500
rect 8800 10400 8900 10500
rect 9000 10400 9100 10500
rect 9200 10400 9300 10500
rect 9400 10400 9500 10500
rect 9600 10400 9700 10500
rect 9800 10400 9900 10500
rect 10000 10400 10100 10500
rect 10200 10400 10300 10500
rect 10400 10400 10500 10500
rect 10600 10400 10700 10500
rect 10800 10400 10900 10500
rect 11000 10400 11100 10500
rect 11200 10400 11300 10500
rect 11400 10400 11500 10500
rect 11600 10400 11700 10500
rect 11800 10400 11900 10500
rect 12000 10400 12100 10500
rect 12200 10400 12300 10500
rect 12400 10400 12500 10500
rect 12600 10400 12700 10500
rect 12800 10400 12900 10500
rect 13000 10400 13100 10500
rect 13200 10400 13300 10500
rect 13400 10400 13500 10500
rect 13600 10400 13700 10500
rect 13800 10400 13900 10500
rect 14000 10400 14100 10500
rect 14200 10400 14300 10500
rect 14400 10400 14500 10500
rect 14600 10400 14700 10500
rect 14800 10400 14900 10500
rect 15000 10400 15100 10500
rect 15200 10400 15300 10500
rect 15400 10400 15500 10500
rect 15600 10400 15700 10500
rect 15800 10400 15900 10500
rect 16000 10400 16100 10500
rect 16200 10400 16300 10500
rect 16400 10400 16500 10500
rect 16600 10400 16700 10500
rect 16800 10400 16900 10500
rect 17000 10400 17100 10500
rect 17200 10400 17300 10500
rect 17400 10400 17500 10500
rect 17600 10400 17700 10500
rect 17800 10400 17900 10500
rect 18000 10400 18100 10500
rect 18200 10400 18300 10500
rect 18400 10400 18500 10500
rect 18600 10400 18700 10500
rect 18800 10400 18900 10500
rect 19000 10400 19100 10500
rect 19200 10400 19300 10500
rect 19400 10400 19500 10500
rect 19600 10400 19700 10500
rect 19800 10400 19900 10500
rect 20000 10400 20100 10500
rect 20200 10400 20300 10500
rect 20400 10400 20500 10500
rect 20600 10400 20700 10500
rect 20800 10400 20900 10500
rect 21000 10400 21100 10500
rect 21200 10400 21300 10500
rect 21400 10400 21500 10500
rect 21600 10400 21700 10500
rect 21800 10400 21900 10500
rect 22000 10400 22100 10500
rect 22200 10400 22300 10500
rect 22400 10400 22500 10500
rect 22600 10400 22700 10500
rect 22800 10400 22900 10500
rect 23000 10400 23100 10500
rect 23200 10400 23300 10500
rect 23400 10400 23500 10500
rect 23600 10400 23700 10500
rect 23800 10400 23900 10500
rect 24000 10400 24100 10500
rect 24200 10400 24300 10500
rect 24400 10400 24500 10500
rect 24600 10400 24700 10500
rect 24800 10400 24900 10500
rect 25000 10400 25100 10500
rect 25200 10400 25300 10500
rect 25400 10400 25500 10500
rect 25600 10400 25700 10500
rect 25800 10400 25900 10500
rect 26000 10400 26100 10500
rect 26200 10400 26300 10500
rect 26400 10400 26500 10500
rect 26600 10400 26700 10500
rect 26800 10400 26900 10500
rect 27000 10400 27100 10500
rect 27200 10400 27300 10500
rect 27400 10400 27500 10500
rect 27600 10400 27700 10500
rect 27800 10400 27900 10500
rect 28000 10400 28100 10500
rect 28200 10400 28300 10500
rect 28400 10400 28500 10500
rect 28600 10400 28700 10500
rect 28800 10400 28900 10500
rect 29000 10400 29100 10500
rect 29200 10400 29300 10500
rect 29400 10400 29500 10500
rect 29600 10400 29700 10500
rect 29800 10400 29900 10500
rect 30000 10400 30100 10500
rect 30200 10400 30300 10500
rect 30400 10400 30500 10500
rect 30600 10400 30700 10500
rect 30800 10400 30900 10500
rect 31000 10400 31100 10500
rect 31200 10400 31300 10500
rect 31400 10400 31500 10500
rect 31600 10400 31700 10500
rect 31800 10400 31900 10500
rect 32000 10400 32100 10500
rect 32200 10400 32300 10500
rect 32400 10400 32500 10500
rect 32600 10400 32700 10500
rect 32800 10400 32900 10500
rect 33000 10400 33100 10500
rect 33200 10400 33324 10500
rect 176 10000 300 10100
rect 400 10000 500 10100
rect 600 10000 700 10100
rect 800 10000 900 10100
rect 1000 10000 1100 10100
rect 1200 10000 1300 10100
rect 1400 10000 1500 10100
rect 1600 10000 1700 10100
rect 1800 10000 1900 10100
rect 2000 10000 2100 10100
rect 2200 10000 2300 10100
rect 2400 10000 2500 10100
rect 2600 10000 2700 10100
rect 2800 10000 2900 10100
rect 3000 10000 3100 10100
rect 3200 10000 3300 10100
rect 3400 10000 3500 10100
rect 3600 10000 3700 10100
rect 3800 10000 3900 10100
rect 4000 10000 4100 10100
rect 4200 10000 4300 10100
rect 4400 10000 4500 10100
rect 4600 10000 4700 10100
rect 4800 10000 4900 10100
rect 5000 10000 5100 10100
rect 5200 10000 5300 10100
rect 5400 10000 5500 10100
rect 5600 10000 5700 10100
rect 5800 10000 5900 10100
rect 6000 10000 6100 10100
rect 6200 10000 6300 10100
rect 6400 10000 6500 10100
rect 6600 10000 6700 10100
rect 6800 10000 6900 10100
rect 7000 10000 7100 10100
rect 7200 10000 7300 10100
rect 7400 10000 7500 10100
rect 7600 10000 7700 10100
rect 7800 10000 7900 10100
rect 8000 10000 8100 10100
rect 8200 10000 8300 10100
rect 8400 10000 8500 10100
rect 8600 10000 8700 10100
rect 8800 10000 8900 10100
rect 9000 10000 9100 10100
rect 9200 10000 9300 10100
rect 9400 10000 9500 10100
rect 9600 10000 9700 10100
rect 9800 10000 9900 10100
rect 10000 10000 10100 10100
rect 10200 10000 10300 10100
rect 10400 10000 10500 10100
rect 10600 10000 10700 10100
rect 10800 10000 10900 10100
rect 11000 10000 11100 10100
rect 11200 10000 11300 10100
rect 11400 10000 11500 10100
rect 11600 10000 11700 10100
rect 11800 10000 11900 10100
rect 12000 10000 12100 10100
rect 12200 10000 12300 10100
rect 12400 10000 12500 10100
rect 12600 10000 12700 10100
rect 12800 10000 12900 10100
rect 13000 10000 13100 10100
rect 13200 10000 13300 10100
rect 13400 10000 13500 10100
rect 13600 10000 13700 10100
rect 13800 10000 13900 10100
rect 14000 10000 14100 10100
rect 14200 10000 14300 10100
rect 14400 10000 14500 10100
rect 14600 10000 14700 10100
rect 14800 10000 14900 10100
rect 15000 10000 15100 10100
rect 15200 10000 15300 10100
rect 15400 10000 15500 10100
rect 15600 10000 15700 10100
rect 15800 10000 15900 10100
rect 16000 10000 16100 10100
rect 16200 10000 16300 10100
rect 16400 10000 16500 10100
rect 16600 10000 16700 10100
rect 16800 10000 16900 10100
rect 17000 10000 17100 10100
rect 17200 10000 17300 10100
rect 17400 10000 17500 10100
rect 17600 10000 17700 10100
rect 17800 10000 17900 10100
rect 18000 10000 18100 10100
rect 18200 10000 18300 10100
rect 18400 10000 18500 10100
rect 18600 10000 18700 10100
rect 18800 10000 18900 10100
rect 19000 10000 19100 10100
rect 19200 10000 19300 10100
rect 19400 10000 19500 10100
rect 19600 10000 19700 10100
rect 19800 10000 19900 10100
rect 20000 10000 20100 10100
rect 20200 10000 20300 10100
rect 20400 10000 20500 10100
rect 20600 10000 20700 10100
rect 20800 10000 20900 10100
rect 21000 10000 21100 10100
rect 21200 10000 21300 10100
rect 21400 10000 21500 10100
rect 21600 10000 21700 10100
rect 21800 10000 21900 10100
rect 22000 10000 22100 10100
rect 22200 10000 22300 10100
rect 22400 10000 22500 10100
rect 22600 10000 22700 10100
rect 22800 10000 22900 10100
rect 23000 10000 23100 10100
rect 23200 10000 23300 10100
rect 23400 10000 23500 10100
rect 23600 10000 23700 10100
rect 23800 10000 23900 10100
rect 24000 10000 24100 10100
rect 24200 10000 24300 10100
rect 24400 10000 24500 10100
rect 24600 10000 24700 10100
rect 24800 10000 24900 10100
rect 25000 10000 25100 10100
rect 25200 10000 25300 10100
rect 25400 10000 25500 10100
rect 25600 10000 25700 10100
rect 25800 10000 25900 10100
rect 26000 10000 26100 10100
rect 26200 10000 26300 10100
rect 26400 10000 26500 10100
rect 26600 10000 26700 10100
rect 26800 10000 26900 10100
rect 27000 10000 27100 10100
rect 27200 10000 27300 10100
rect 27400 10000 27500 10100
rect 27600 10000 27700 10100
rect 27800 10000 27900 10100
rect 28000 10000 28100 10100
rect 28200 10000 28300 10100
rect 28400 10000 28500 10100
rect 28600 10000 28700 10100
rect 28800 10000 28900 10100
rect 29000 10000 29100 10100
rect 29200 10000 29300 10100
rect 29400 10000 29500 10100
rect 29600 10000 29700 10100
rect 29800 10000 29900 10100
rect 30000 10000 30100 10100
rect 30200 10000 30300 10100
rect 30400 10000 30500 10100
rect 30600 10000 30700 10100
rect 30800 10000 30900 10100
rect 31000 10000 31100 10100
rect 31200 10000 31300 10100
rect 31400 10000 31500 10100
rect 31600 10000 31700 10100
rect 31800 10000 31900 10100
rect 32000 10000 32100 10100
rect 32200 10000 32300 10100
rect 32400 10000 32500 10100
rect 32600 10000 32700 10100
rect 32800 10000 32900 10100
rect 33000 10000 33100 10100
rect 33200 10000 33300 10100
rect 33400 10000 33500 10100
rect 33600 10000 33700 10100
rect 33800 10000 33900 10100
rect 34000 10000 34100 10100
rect 34200 10000 34300 10100
rect 34400 10000 34500 10100
rect 34600 10000 34700 10100
rect 34800 10000 34900 10100
rect 35000 10000 35100 10100
rect 35200 10000 35300 10100
rect 35400 10000 35500 10100
rect 35600 10000 35700 10100
rect 35800 10000 35900 10100
rect 36000 10000 36124 10100
rect 200 9900 300 10000
rect 200 9700 300 9800
rect 200 9500 300 9600
rect 200 9300 300 9400
rect 200 9100 300 9200
rect 200 8900 300 9000
rect 200 8700 300 8800
rect 200 8500 300 8600
rect 200 8300 300 8400
rect 200 8100 300 8200
rect 200 7900 300 8000
rect 200 7700 300 7800
rect 200 7500 300 7600
rect 200 7300 300 7400
rect 200 7100 300 7200
rect 200 6900 300 7000
rect 200 6700 300 6800
rect 200 6500 300 6600
rect 200 6300 300 6400
rect 200 6100 300 6200
rect 36000 9900 36100 10000
rect 36000 9700 36100 9800
rect 36000 9500 36100 9600
rect 36000 9300 36100 9400
rect 36000 9100 36100 9200
rect 36000 8900 36100 9000
rect 36000 8700 36100 8800
rect 36000 8500 36100 8600
rect 36000 8300 36100 8400
rect 36000 8100 36100 8200
rect 36000 7900 36100 8000
rect 36000 7700 36100 7800
rect 36000 7500 36100 7600
rect 36000 7300 36100 7400
rect 36000 7100 36100 7200
rect 36000 6900 36100 7000
rect 36000 6700 36100 6800
rect 36000 6500 36100 6600
rect 36000 6300 36100 6400
rect 36000 6100 36100 6200
rect 176 6000 300 6100
rect 400 6000 500 6100
rect 600 6000 700 6100
rect 800 6000 900 6100
rect 1000 6000 1100 6100
rect 1200 6000 1300 6100
rect 1400 6000 1500 6100
rect 1600 6000 1700 6100
rect 1800 6000 1900 6100
rect 2000 6000 2100 6100
rect 2200 6000 2300 6100
rect 2400 6000 2500 6100
rect 2600 6000 2700 6100
rect 2800 6000 2900 6100
rect 3000 6000 3100 6100
rect 3200 6000 3300 6100
rect 3400 6000 3500 6100
rect 3600 6000 3700 6100
rect 3800 6000 3900 6100
rect 4000 6000 4100 6100
rect 4200 6000 4300 6100
rect 4400 6000 4500 6100
rect 4600 6000 4700 6100
rect 4800 6000 4900 6100
rect 5000 6000 5100 6100
rect 5200 6000 5300 6100
rect 5400 6000 5500 6100
rect 5600 6000 5700 6100
rect 5800 6000 5900 6100
rect 6000 6000 6100 6100
rect 6200 6000 6300 6100
rect 6400 6000 6500 6100
rect 6600 6000 6700 6100
rect 6800 6000 6900 6100
rect 7000 6000 7100 6100
rect 7200 6000 7300 6100
rect 7400 6000 7500 6100
rect 7600 6000 7700 6100
rect 7800 6000 7900 6100
rect 8000 6000 8100 6100
rect 8200 6000 8300 6100
rect 8400 6000 8500 6100
rect 8600 6000 8700 6100
rect 8800 6000 8900 6100
rect 9000 6000 9100 6100
rect 9200 6000 9300 6100
rect 9400 6000 9500 6100
rect 9600 6000 9700 6100
rect 9800 6000 9900 6100
rect 10000 6000 10100 6100
rect 10200 6000 10300 6100
rect 10400 6000 10500 6100
rect 10600 6000 10700 6100
rect 10800 6000 10900 6100
rect 11000 6000 11100 6100
rect 11200 6000 11300 6100
rect 11400 6000 11500 6100
rect 11600 6000 11700 6100
rect 11800 6000 11900 6100
rect 12000 6000 12100 6100
rect 12200 6000 12300 6100
rect 12400 6000 12500 6100
rect 12600 6000 12700 6100
rect 12800 6000 12900 6100
rect 13000 6000 13100 6100
rect 13200 6000 13300 6100
rect 13400 6000 13500 6100
rect 13600 6000 13700 6100
rect 13800 6000 13900 6100
rect 14000 6000 14100 6100
rect 14200 6000 14300 6100
rect 14400 6000 14500 6100
rect 14600 6000 14700 6100
rect 14800 6000 14900 6100
rect 15000 6000 15100 6100
rect 15200 6000 15300 6100
rect 15400 6000 15500 6100
rect 15600 6000 15700 6100
rect 15800 6000 15900 6100
rect 16000 6000 16100 6100
rect 16200 6000 16300 6100
rect 16400 6000 16500 6100
rect 16600 6000 16700 6100
rect 16800 6000 16900 6100
rect 17000 6000 17100 6100
rect 17200 6000 17300 6100
rect 17400 6000 17500 6100
rect 17600 6000 17700 6100
rect 17800 6000 17900 6100
rect 18000 6000 18100 6100
rect 18200 6000 18300 6100
rect 18400 6000 18500 6100
rect 18600 6000 18700 6100
rect 18800 6000 18900 6100
rect 19000 6000 19100 6100
rect 19200 6000 19300 6100
rect 19400 6000 19500 6100
rect 19600 6000 19700 6100
rect 19800 6000 19900 6100
rect 20000 6000 20100 6100
rect 20200 6000 20300 6100
rect 20400 6000 20500 6100
rect 20600 6000 20700 6100
rect 20800 6000 20900 6100
rect 21000 6000 21100 6100
rect 21200 6000 21300 6100
rect 21400 6000 21500 6100
rect 21600 6000 21700 6100
rect 21800 6000 21900 6100
rect 22000 6000 22100 6100
rect 22200 6000 22300 6100
rect 22400 6000 22500 6100
rect 22600 6000 22700 6100
rect 22800 6000 22900 6100
rect 23000 6000 23100 6100
rect 23200 6000 23300 6100
rect 23400 6000 23500 6100
rect 23600 6000 23700 6100
rect 23800 6000 23900 6100
rect 24000 6000 24100 6100
rect 24200 6000 24300 6100
rect 24400 6000 24500 6100
rect 24600 6000 24700 6100
rect 24800 6000 24900 6100
rect 25000 6000 25100 6100
rect 25200 6000 25300 6100
rect 25400 6000 25500 6100
rect 25600 6000 25700 6100
rect 25800 6000 25900 6100
rect 26000 6000 26100 6100
rect 26200 6000 26300 6100
rect 26400 6000 26500 6100
rect 26600 6000 26700 6100
rect 26800 6000 26900 6100
rect 27000 6000 27100 6100
rect 27200 6000 27300 6100
rect 27400 6000 27500 6100
rect 27600 6000 27700 6100
rect 27800 6000 27900 6100
rect 28000 6000 28100 6100
rect 28200 6000 28300 6100
rect 28400 6000 28500 6100
rect 28600 6000 28700 6100
rect 28800 6000 28900 6100
rect 29000 6000 29100 6100
rect 29200 6000 29300 6100
rect 29400 6000 29500 6100
rect 29600 6000 29700 6100
rect 29800 6000 29900 6100
rect 30000 6000 30100 6100
rect 30200 6000 30300 6100
rect 30400 6000 30500 6100
rect 30600 6000 30700 6100
rect 30800 6000 30900 6100
rect 31000 6000 31100 6100
rect 31200 6000 31300 6100
rect 31400 6000 31500 6100
rect 31600 6000 31700 6100
rect 31800 6000 31900 6100
rect 32000 6000 32100 6100
rect 32200 6000 32300 6100
rect 32400 6000 32500 6100
rect 32600 6000 32700 6100
rect 32800 6000 32900 6100
rect 33000 6000 33100 6100
rect 33200 6000 33300 6100
rect 33400 6000 33500 6100
rect 33600 6000 33700 6100
rect 33800 6000 33900 6100
rect 34000 6000 34100 6100
rect 34200 6000 34300 6100
rect 34400 6000 34500 6100
rect 34600 6000 34700 6100
rect 34800 6000 34900 6100
rect 35000 6000 35100 6100
rect 35200 6000 35300 6100
rect 35400 6000 35500 6100
rect 35600 6000 35700 6100
rect 35800 6000 35900 6100
rect 36000 6000 36124 6100
<< psubdiffcont >>
rect 3300 14400 3400 14500
rect 3500 14400 3600 14500
rect 3700 14400 3800 14500
rect 3900 14400 4000 14500
rect 4100 14400 4200 14500
rect 4300 14400 4400 14500
rect 4500 14400 4600 14500
rect 4700 14400 4800 14500
rect 4900 14400 5000 14500
rect 5100 14400 5200 14500
rect 5300 14400 5400 14500
rect 5500 14400 5600 14500
rect 5700 14400 5800 14500
rect 5900 14400 6000 14500
rect 6100 14400 6200 14500
rect 6300 14400 6400 14500
rect 6500 14400 6600 14500
rect 6700 14400 6800 14500
rect 6900 14400 7000 14500
rect 7100 14400 7200 14500
rect 7300 14400 7400 14500
rect 7500 14400 7600 14500
rect 7700 14400 7800 14500
rect 7900 14400 8000 14500
rect 8100 14400 8200 14500
rect 8300 14400 8400 14500
rect 8500 14400 8600 14500
rect 8700 14400 8800 14500
rect 8900 14400 9000 14500
rect 9100 14400 9200 14500
rect 9300 14400 9400 14500
rect 9500 14400 9600 14500
rect 9700 14400 9800 14500
rect 9900 14400 10000 14500
rect 10100 14400 10200 14500
rect 10300 14400 10400 14500
rect 10500 14400 10600 14500
rect 10700 14400 10800 14500
rect 10900 14400 11000 14500
rect 11100 14400 11200 14500
rect 11300 14400 11400 14500
rect 11500 14400 11600 14500
rect 11700 14400 11800 14500
rect 11900 14400 12000 14500
rect 12100 14400 12200 14500
rect 12300 14400 12400 14500
rect 12500 14400 12600 14500
rect 12700 14400 12800 14500
rect 12900 14400 13000 14500
rect 13100 14400 13200 14500
rect 13300 14400 13400 14500
rect 13500 14400 13600 14500
rect 13700 14400 13800 14500
rect 13900 14400 14000 14500
rect 14100 14400 14200 14500
rect 14300 14400 14400 14500
rect 14500 14400 14600 14500
rect 14700 14400 14800 14500
rect 14900 14400 15000 14500
rect 15100 14400 15200 14500
rect 15300 14400 15400 14500
rect 15500 14400 15600 14500
rect 15700 14400 15800 14500
rect 15900 14400 16000 14500
rect 16100 14400 16200 14500
rect 16300 14400 16400 14500
rect 16500 14400 16600 14500
rect 16700 14400 16800 14500
rect 16900 14400 17000 14500
rect 17100 14400 17200 14500
rect 17300 14400 17400 14500
rect 17500 14400 17600 14500
rect 17700 14400 17800 14500
rect 17900 14400 18000 14500
rect 18100 14400 18200 14500
rect 18300 14400 18400 14500
rect 18500 14400 18600 14500
rect 18700 14400 18800 14500
rect 18900 14400 19000 14500
rect 19100 14400 19200 14500
rect 19300 14400 19400 14500
rect 19500 14400 19600 14500
rect 19700 14400 19800 14500
rect 19900 14400 20000 14500
rect 20100 14400 20200 14500
rect 20300 14400 20400 14500
rect 20500 14400 20600 14500
rect 20700 14400 20800 14500
rect 20900 14400 21000 14500
rect 21100 14400 21200 14500
rect 21300 14400 21400 14500
rect 21500 14400 21600 14500
rect 21700 14400 21800 14500
rect 21900 14400 22000 14500
rect 22100 14400 22200 14500
rect 22300 14400 22400 14500
rect 22500 14400 22600 14500
rect 22700 14400 22800 14500
rect 22900 14400 23000 14500
rect 23100 14400 23200 14500
rect 23300 14400 23400 14500
rect 23500 14400 23600 14500
rect 23700 14400 23800 14500
rect 23900 14400 24000 14500
rect 24100 14400 24200 14500
rect 24300 14400 24400 14500
rect 24500 14400 24600 14500
rect 24700 14400 24800 14500
rect 24900 14400 25000 14500
rect 25100 14400 25200 14500
rect 25300 14400 25400 14500
rect 25500 14400 25600 14500
rect 25700 14400 25800 14500
rect 25900 14400 26000 14500
rect 26100 14400 26200 14500
rect 26300 14400 26400 14500
rect 26500 14400 26600 14500
rect 26700 14400 26800 14500
rect 26900 14400 27000 14500
rect 27100 14400 27200 14500
rect 27300 14400 27400 14500
rect 27500 14400 27600 14500
rect 27700 14400 27800 14500
rect 27900 14400 28000 14500
rect 28100 14400 28200 14500
rect 28300 14400 28400 14500
rect 28500 14400 28600 14500
rect 28700 14400 28800 14500
rect 28900 14400 29000 14500
rect 29100 14400 29200 14500
rect 29300 14400 29400 14500
rect 29500 14400 29600 14500
rect 29700 14400 29800 14500
rect 29900 14400 30000 14500
rect 30100 14400 30200 14500
rect 30300 14400 30400 14500
rect 30500 14400 30600 14500
rect 30700 14400 30800 14500
rect 30900 14400 31000 14500
rect 31100 14400 31200 14500
rect 31300 14400 31400 14500
rect 31500 14400 31600 14500
rect 31700 14400 31800 14500
rect 31900 14400 32000 14500
rect 32100 14400 32200 14500
rect 32300 14400 32400 14500
rect 32500 14400 32600 14500
rect 32700 14400 32800 14500
rect 32900 14400 33000 14500
rect 33100 14400 33200 14500
rect 3200 14200 3300 14300
rect 3200 14000 3300 14100
rect 3200 13800 3300 13900
rect 3200 13600 3300 13700
rect 3200 13400 3300 13500
rect 3200 13200 3300 13300
rect 3200 13000 3300 13100
rect 3200 12800 3300 12900
rect 3200 12600 3300 12700
rect 3200 12400 3300 12500
rect 3200 12200 3300 12300
rect 3200 12000 3300 12100
rect 3200 11800 3300 11900
rect 3200 11600 3300 11700
rect 3200 11400 3300 11500
rect 3200 11200 3300 11300
rect 3200 11000 3300 11100
rect 3200 10800 3300 10900
rect 3200 10600 3300 10700
rect 33200 14200 33300 14300
rect 33200 14000 33300 14100
rect 33200 13800 33300 13900
rect 33200 13600 33300 13700
rect 33200 13400 33300 13500
rect 33200 13200 33300 13300
rect 33200 13000 33300 13100
rect 33200 12800 33300 12900
rect 33200 12600 33300 12700
rect 33200 12400 33300 12500
rect 33200 12200 33300 12300
rect 33200 12000 33300 12100
rect 33200 11800 33300 11900
rect 33200 11600 33300 11700
rect 33200 11400 33300 11500
rect 33200 11200 33300 11300
rect 33200 11000 33300 11100
rect 33200 10800 33300 10900
rect 33200 10600 33300 10700
rect 3300 10400 3400 10500
rect 3500 10400 3600 10500
rect 3700 10400 3800 10500
rect 3900 10400 4000 10500
rect 4100 10400 4200 10500
rect 4300 10400 4400 10500
rect 4500 10400 4600 10500
rect 4700 10400 4800 10500
rect 4900 10400 5000 10500
rect 5100 10400 5200 10500
rect 5300 10400 5400 10500
rect 5500 10400 5600 10500
rect 5700 10400 5800 10500
rect 5900 10400 6000 10500
rect 6100 10400 6200 10500
rect 6300 10400 6400 10500
rect 6500 10400 6600 10500
rect 6700 10400 6800 10500
rect 6900 10400 7000 10500
rect 7100 10400 7200 10500
rect 7300 10400 7400 10500
rect 7500 10400 7600 10500
rect 7700 10400 7800 10500
rect 7900 10400 8000 10500
rect 8100 10400 8200 10500
rect 8300 10400 8400 10500
rect 8500 10400 8600 10500
rect 8700 10400 8800 10500
rect 8900 10400 9000 10500
rect 9100 10400 9200 10500
rect 9300 10400 9400 10500
rect 9500 10400 9600 10500
rect 9700 10400 9800 10500
rect 9900 10400 10000 10500
rect 10100 10400 10200 10500
rect 10300 10400 10400 10500
rect 10500 10400 10600 10500
rect 10700 10400 10800 10500
rect 10900 10400 11000 10500
rect 11100 10400 11200 10500
rect 11300 10400 11400 10500
rect 11500 10400 11600 10500
rect 11700 10400 11800 10500
rect 11900 10400 12000 10500
rect 12100 10400 12200 10500
rect 12300 10400 12400 10500
rect 12500 10400 12600 10500
rect 12700 10400 12800 10500
rect 12900 10400 13000 10500
rect 13100 10400 13200 10500
rect 13300 10400 13400 10500
rect 13500 10400 13600 10500
rect 13700 10400 13800 10500
rect 13900 10400 14000 10500
rect 14100 10400 14200 10500
rect 14300 10400 14400 10500
rect 14500 10400 14600 10500
rect 14700 10400 14800 10500
rect 14900 10400 15000 10500
rect 15100 10400 15200 10500
rect 15300 10400 15400 10500
rect 15500 10400 15600 10500
rect 15700 10400 15800 10500
rect 15900 10400 16000 10500
rect 16100 10400 16200 10500
rect 16300 10400 16400 10500
rect 16500 10400 16600 10500
rect 16700 10400 16800 10500
rect 16900 10400 17000 10500
rect 17100 10400 17200 10500
rect 17300 10400 17400 10500
rect 17500 10400 17600 10500
rect 17700 10400 17800 10500
rect 17900 10400 18000 10500
rect 18100 10400 18200 10500
rect 18300 10400 18400 10500
rect 18500 10400 18600 10500
rect 18700 10400 18800 10500
rect 18900 10400 19000 10500
rect 19100 10400 19200 10500
rect 19300 10400 19400 10500
rect 19500 10400 19600 10500
rect 19700 10400 19800 10500
rect 19900 10400 20000 10500
rect 20100 10400 20200 10500
rect 20300 10400 20400 10500
rect 20500 10400 20600 10500
rect 20700 10400 20800 10500
rect 20900 10400 21000 10500
rect 21100 10400 21200 10500
rect 21300 10400 21400 10500
rect 21500 10400 21600 10500
rect 21700 10400 21800 10500
rect 21900 10400 22000 10500
rect 22100 10400 22200 10500
rect 22300 10400 22400 10500
rect 22500 10400 22600 10500
rect 22700 10400 22800 10500
rect 22900 10400 23000 10500
rect 23100 10400 23200 10500
rect 23300 10400 23400 10500
rect 23500 10400 23600 10500
rect 23700 10400 23800 10500
rect 23900 10400 24000 10500
rect 24100 10400 24200 10500
rect 24300 10400 24400 10500
rect 24500 10400 24600 10500
rect 24700 10400 24800 10500
rect 24900 10400 25000 10500
rect 25100 10400 25200 10500
rect 25300 10400 25400 10500
rect 25500 10400 25600 10500
rect 25700 10400 25800 10500
rect 25900 10400 26000 10500
rect 26100 10400 26200 10500
rect 26300 10400 26400 10500
rect 26500 10400 26600 10500
rect 26700 10400 26800 10500
rect 26900 10400 27000 10500
rect 27100 10400 27200 10500
rect 27300 10400 27400 10500
rect 27500 10400 27600 10500
rect 27700 10400 27800 10500
rect 27900 10400 28000 10500
rect 28100 10400 28200 10500
rect 28300 10400 28400 10500
rect 28500 10400 28600 10500
rect 28700 10400 28800 10500
rect 28900 10400 29000 10500
rect 29100 10400 29200 10500
rect 29300 10400 29400 10500
rect 29500 10400 29600 10500
rect 29700 10400 29800 10500
rect 29900 10400 30000 10500
rect 30100 10400 30200 10500
rect 30300 10400 30400 10500
rect 30500 10400 30600 10500
rect 30700 10400 30800 10500
rect 30900 10400 31000 10500
rect 31100 10400 31200 10500
rect 31300 10400 31400 10500
rect 31500 10400 31600 10500
rect 31700 10400 31800 10500
rect 31900 10400 32000 10500
rect 32100 10400 32200 10500
rect 32300 10400 32400 10500
rect 32500 10400 32600 10500
rect 32700 10400 32800 10500
rect 32900 10400 33000 10500
rect 33100 10400 33200 10500
rect 300 10000 400 10100
rect 500 10000 600 10100
rect 700 10000 800 10100
rect 900 10000 1000 10100
rect 1100 10000 1200 10100
rect 1300 10000 1400 10100
rect 1500 10000 1600 10100
rect 1700 10000 1800 10100
rect 1900 10000 2000 10100
rect 2100 10000 2200 10100
rect 2300 10000 2400 10100
rect 2500 10000 2600 10100
rect 2700 10000 2800 10100
rect 2900 10000 3000 10100
rect 3100 10000 3200 10100
rect 3300 10000 3400 10100
rect 3500 10000 3600 10100
rect 3700 10000 3800 10100
rect 3900 10000 4000 10100
rect 4100 10000 4200 10100
rect 4300 10000 4400 10100
rect 4500 10000 4600 10100
rect 4700 10000 4800 10100
rect 4900 10000 5000 10100
rect 5100 10000 5200 10100
rect 5300 10000 5400 10100
rect 5500 10000 5600 10100
rect 5700 10000 5800 10100
rect 5900 10000 6000 10100
rect 6100 10000 6200 10100
rect 6300 10000 6400 10100
rect 6500 10000 6600 10100
rect 6700 10000 6800 10100
rect 6900 10000 7000 10100
rect 7100 10000 7200 10100
rect 7300 10000 7400 10100
rect 7500 10000 7600 10100
rect 7700 10000 7800 10100
rect 7900 10000 8000 10100
rect 8100 10000 8200 10100
rect 8300 10000 8400 10100
rect 8500 10000 8600 10100
rect 8700 10000 8800 10100
rect 8900 10000 9000 10100
rect 9100 10000 9200 10100
rect 9300 10000 9400 10100
rect 9500 10000 9600 10100
rect 9700 10000 9800 10100
rect 9900 10000 10000 10100
rect 10100 10000 10200 10100
rect 10300 10000 10400 10100
rect 10500 10000 10600 10100
rect 10700 10000 10800 10100
rect 10900 10000 11000 10100
rect 11100 10000 11200 10100
rect 11300 10000 11400 10100
rect 11500 10000 11600 10100
rect 11700 10000 11800 10100
rect 11900 10000 12000 10100
rect 12100 10000 12200 10100
rect 12300 10000 12400 10100
rect 12500 10000 12600 10100
rect 12700 10000 12800 10100
rect 12900 10000 13000 10100
rect 13100 10000 13200 10100
rect 13300 10000 13400 10100
rect 13500 10000 13600 10100
rect 13700 10000 13800 10100
rect 13900 10000 14000 10100
rect 14100 10000 14200 10100
rect 14300 10000 14400 10100
rect 14500 10000 14600 10100
rect 14700 10000 14800 10100
rect 14900 10000 15000 10100
rect 15100 10000 15200 10100
rect 15300 10000 15400 10100
rect 15500 10000 15600 10100
rect 15700 10000 15800 10100
rect 15900 10000 16000 10100
rect 16100 10000 16200 10100
rect 16300 10000 16400 10100
rect 16500 10000 16600 10100
rect 16700 10000 16800 10100
rect 16900 10000 17000 10100
rect 17100 10000 17200 10100
rect 17300 10000 17400 10100
rect 17500 10000 17600 10100
rect 17700 10000 17800 10100
rect 17900 10000 18000 10100
rect 18100 10000 18200 10100
rect 18300 10000 18400 10100
rect 18500 10000 18600 10100
rect 18700 10000 18800 10100
rect 18900 10000 19000 10100
rect 19100 10000 19200 10100
rect 19300 10000 19400 10100
rect 19500 10000 19600 10100
rect 19700 10000 19800 10100
rect 19900 10000 20000 10100
rect 20100 10000 20200 10100
rect 20300 10000 20400 10100
rect 20500 10000 20600 10100
rect 20700 10000 20800 10100
rect 20900 10000 21000 10100
rect 21100 10000 21200 10100
rect 21300 10000 21400 10100
rect 21500 10000 21600 10100
rect 21700 10000 21800 10100
rect 21900 10000 22000 10100
rect 22100 10000 22200 10100
rect 22300 10000 22400 10100
rect 22500 10000 22600 10100
rect 22700 10000 22800 10100
rect 22900 10000 23000 10100
rect 23100 10000 23200 10100
rect 23300 10000 23400 10100
rect 23500 10000 23600 10100
rect 23700 10000 23800 10100
rect 23900 10000 24000 10100
rect 24100 10000 24200 10100
rect 24300 10000 24400 10100
rect 24500 10000 24600 10100
rect 24700 10000 24800 10100
rect 24900 10000 25000 10100
rect 25100 10000 25200 10100
rect 25300 10000 25400 10100
rect 25500 10000 25600 10100
rect 25700 10000 25800 10100
rect 25900 10000 26000 10100
rect 26100 10000 26200 10100
rect 26300 10000 26400 10100
rect 26500 10000 26600 10100
rect 26700 10000 26800 10100
rect 26900 10000 27000 10100
rect 27100 10000 27200 10100
rect 27300 10000 27400 10100
rect 27500 10000 27600 10100
rect 27700 10000 27800 10100
rect 27900 10000 28000 10100
rect 28100 10000 28200 10100
rect 28300 10000 28400 10100
rect 28500 10000 28600 10100
rect 28700 10000 28800 10100
rect 28900 10000 29000 10100
rect 29100 10000 29200 10100
rect 29300 10000 29400 10100
rect 29500 10000 29600 10100
rect 29700 10000 29800 10100
rect 29900 10000 30000 10100
rect 30100 10000 30200 10100
rect 30300 10000 30400 10100
rect 30500 10000 30600 10100
rect 30700 10000 30800 10100
rect 30900 10000 31000 10100
rect 31100 10000 31200 10100
rect 31300 10000 31400 10100
rect 31500 10000 31600 10100
rect 31700 10000 31800 10100
rect 31900 10000 32000 10100
rect 32100 10000 32200 10100
rect 32300 10000 32400 10100
rect 32500 10000 32600 10100
rect 32700 10000 32800 10100
rect 32900 10000 33000 10100
rect 33100 10000 33200 10100
rect 33300 10000 33400 10100
rect 33500 10000 33600 10100
rect 33700 10000 33800 10100
rect 33900 10000 34000 10100
rect 34100 10000 34200 10100
rect 34300 10000 34400 10100
rect 34500 10000 34600 10100
rect 34700 10000 34800 10100
rect 34900 10000 35000 10100
rect 35100 10000 35200 10100
rect 35300 10000 35400 10100
rect 35500 10000 35600 10100
rect 35700 10000 35800 10100
rect 35900 10000 36000 10100
rect 200 9800 300 9900
rect 200 9600 300 9700
rect 200 9400 300 9500
rect 200 9200 300 9300
rect 200 9000 300 9100
rect 200 8800 300 8900
rect 200 8600 300 8700
rect 200 8400 300 8500
rect 200 8200 300 8300
rect 200 8000 300 8100
rect 200 7800 300 7900
rect 200 7600 300 7700
rect 200 7400 300 7500
rect 200 7200 300 7300
rect 200 7000 300 7100
rect 200 6800 300 6900
rect 200 6600 300 6700
rect 200 6400 300 6500
rect 200 6200 300 6300
rect 36000 9800 36100 9900
rect 36000 9600 36100 9700
rect 36000 9400 36100 9500
rect 36000 9200 36100 9300
rect 36000 9000 36100 9100
rect 36000 8800 36100 8900
rect 36000 8600 36100 8700
rect 36000 8400 36100 8500
rect 36000 8200 36100 8300
rect 36000 8000 36100 8100
rect 36000 7800 36100 7900
rect 36000 7600 36100 7700
rect 36000 7400 36100 7500
rect 36000 7200 36100 7300
rect 36000 7000 36100 7100
rect 36000 6800 36100 6900
rect 36000 6600 36100 6700
rect 36000 6400 36100 6500
rect 36000 6200 36100 6300
rect 300 6000 400 6100
rect 500 6000 600 6100
rect 700 6000 800 6100
rect 900 6000 1000 6100
rect 1100 6000 1200 6100
rect 1300 6000 1400 6100
rect 1500 6000 1600 6100
rect 1700 6000 1800 6100
rect 1900 6000 2000 6100
rect 2100 6000 2200 6100
rect 2300 6000 2400 6100
rect 2500 6000 2600 6100
rect 2700 6000 2800 6100
rect 2900 6000 3000 6100
rect 3100 6000 3200 6100
rect 3300 6000 3400 6100
rect 3500 6000 3600 6100
rect 3700 6000 3800 6100
rect 3900 6000 4000 6100
rect 4100 6000 4200 6100
rect 4300 6000 4400 6100
rect 4500 6000 4600 6100
rect 4700 6000 4800 6100
rect 4900 6000 5000 6100
rect 5100 6000 5200 6100
rect 5300 6000 5400 6100
rect 5500 6000 5600 6100
rect 5700 6000 5800 6100
rect 5900 6000 6000 6100
rect 6100 6000 6200 6100
rect 6300 6000 6400 6100
rect 6500 6000 6600 6100
rect 6700 6000 6800 6100
rect 6900 6000 7000 6100
rect 7100 6000 7200 6100
rect 7300 6000 7400 6100
rect 7500 6000 7600 6100
rect 7700 6000 7800 6100
rect 7900 6000 8000 6100
rect 8100 6000 8200 6100
rect 8300 6000 8400 6100
rect 8500 6000 8600 6100
rect 8700 6000 8800 6100
rect 8900 6000 9000 6100
rect 9100 6000 9200 6100
rect 9300 6000 9400 6100
rect 9500 6000 9600 6100
rect 9700 6000 9800 6100
rect 9900 6000 10000 6100
rect 10100 6000 10200 6100
rect 10300 6000 10400 6100
rect 10500 6000 10600 6100
rect 10700 6000 10800 6100
rect 10900 6000 11000 6100
rect 11100 6000 11200 6100
rect 11300 6000 11400 6100
rect 11500 6000 11600 6100
rect 11700 6000 11800 6100
rect 11900 6000 12000 6100
rect 12100 6000 12200 6100
rect 12300 6000 12400 6100
rect 12500 6000 12600 6100
rect 12700 6000 12800 6100
rect 12900 6000 13000 6100
rect 13100 6000 13200 6100
rect 13300 6000 13400 6100
rect 13500 6000 13600 6100
rect 13700 6000 13800 6100
rect 13900 6000 14000 6100
rect 14100 6000 14200 6100
rect 14300 6000 14400 6100
rect 14500 6000 14600 6100
rect 14700 6000 14800 6100
rect 14900 6000 15000 6100
rect 15100 6000 15200 6100
rect 15300 6000 15400 6100
rect 15500 6000 15600 6100
rect 15700 6000 15800 6100
rect 15900 6000 16000 6100
rect 16100 6000 16200 6100
rect 16300 6000 16400 6100
rect 16500 6000 16600 6100
rect 16700 6000 16800 6100
rect 16900 6000 17000 6100
rect 17100 6000 17200 6100
rect 17300 6000 17400 6100
rect 17500 6000 17600 6100
rect 17700 6000 17800 6100
rect 17900 6000 18000 6100
rect 18100 6000 18200 6100
rect 18300 6000 18400 6100
rect 18500 6000 18600 6100
rect 18700 6000 18800 6100
rect 18900 6000 19000 6100
rect 19100 6000 19200 6100
rect 19300 6000 19400 6100
rect 19500 6000 19600 6100
rect 19700 6000 19800 6100
rect 19900 6000 20000 6100
rect 20100 6000 20200 6100
rect 20300 6000 20400 6100
rect 20500 6000 20600 6100
rect 20700 6000 20800 6100
rect 20900 6000 21000 6100
rect 21100 6000 21200 6100
rect 21300 6000 21400 6100
rect 21500 6000 21600 6100
rect 21700 6000 21800 6100
rect 21900 6000 22000 6100
rect 22100 6000 22200 6100
rect 22300 6000 22400 6100
rect 22500 6000 22600 6100
rect 22700 6000 22800 6100
rect 22900 6000 23000 6100
rect 23100 6000 23200 6100
rect 23300 6000 23400 6100
rect 23500 6000 23600 6100
rect 23700 6000 23800 6100
rect 23900 6000 24000 6100
rect 24100 6000 24200 6100
rect 24300 6000 24400 6100
rect 24500 6000 24600 6100
rect 24700 6000 24800 6100
rect 24900 6000 25000 6100
rect 25100 6000 25200 6100
rect 25300 6000 25400 6100
rect 25500 6000 25600 6100
rect 25700 6000 25800 6100
rect 25900 6000 26000 6100
rect 26100 6000 26200 6100
rect 26300 6000 26400 6100
rect 26500 6000 26600 6100
rect 26700 6000 26800 6100
rect 26900 6000 27000 6100
rect 27100 6000 27200 6100
rect 27300 6000 27400 6100
rect 27500 6000 27600 6100
rect 27700 6000 27800 6100
rect 27900 6000 28000 6100
rect 28100 6000 28200 6100
rect 28300 6000 28400 6100
rect 28500 6000 28600 6100
rect 28700 6000 28800 6100
rect 28900 6000 29000 6100
rect 29100 6000 29200 6100
rect 29300 6000 29400 6100
rect 29500 6000 29600 6100
rect 29700 6000 29800 6100
rect 29900 6000 30000 6100
rect 30100 6000 30200 6100
rect 30300 6000 30400 6100
rect 30500 6000 30600 6100
rect 30700 6000 30800 6100
rect 30900 6000 31000 6100
rect 31100 6000 31200 6100
rect 31300 6000 31400 6100
rect 31500 6000 31600 6100
rect 31700 6000 31800 6100
rect 31900 6000 32000 6100
rect 32100 6000 32200 6100
rect 32300 6000 32400 6100
rect 32500 6000 32600 6100
rect 32700 6000 32800 6100
rect 32900 6000 33000 6100
rect 33100 6000 33200 6100
rect 33300 6000 33400 6100
rect 33500 6000 33600 6100
rect 33700 6000 33800 6100
rect 33900 6000 34000 6100
rect 34100 6000 34200 6100
rect 34300 6000 34400 6100
rect 34500 6000 34600 6100
rect 34700 6000 34800 6100
rect 34900 6000 35000 6100
rect 35100 6000 35200 6100
rect 35300 6000 35400 6100
rect 35500 6000 35600 6100
rect 35700 6000 35800 6100
rect 35900 6000 36000 6100
<< locali >>
rect 3184 14400 3300 14500
rect 3400 14400 3500 14500
rect 3600 14400 3700 14500
rect 3800 14400 3900 14500
rect 4000 14400 4100 14500
rect 4200 14400 4300 14500
rect 4400 14400 4500 14500
rect 4600 14400 4700 14500
rect 4800 14400 4900 14500
rect 5000 14400 5100 14500
rect 5200 14400 5300 14500
rect 5400 14400 5500 14500
rect 5600 14400 5700 14500
rect 5800 14400 5900 14500
rect 6000 14400 6100 14500
rect 6200 14400 6300 14500
rect 6400 14400 6500 14500
rect 6600 14400 6700 14500
rect 6800 14400 6900 14500
rect 7000 14400 7100 14500
rect 7200 14400 7300 14500
rect 7400 14400 7500 14500
rect 7600 14400 7700 14500
rect 7800 14400 7900 14500
rect 8000 14400 8100 14500
rect 8200 14400 8300 14500
rect 8400 14400 8500 14500
rect 8600 14400 8700 14500
rect 8800 14400 8900 14500
rect 9000 14400 9100 14500
rect 9200 14400 9300 14500
rect 9400 14400 9500 14500
rect 9600 14400 9700 14500
rect 9800 14400 9900 14500
rect 10000 14400 10100 14500
rect 10200 14400 10300 14500
rect 10400 14400 10500 14500
rect 10600 14400 10700 14500
rect 10800 14400 10900 14500
rect 11000 14400 11100 14500
rect 11200 14400 11300 14500
rect 11400 14400 11500 14500
rect 11600 14400 11700 14500
rect 11800 14400 11900 14500
rect 12000 14400 12100 14500
rect 12200 14400 12300 14500
rect 12400 14400 12500 14500
rect 12600 14400 12700 14500
rect 12800 14400 12900 14500
rect 13000 14400 13100 14500
rect 13200 14400 13300 14500
rect 13400 14400 13500 14500
rect 13600 14400 13700 14500
rect 13800 14400 13900 14500
rect 14000 14400 14100 14500
rect 14200 14400 14300 14500
rect 14400 14400 14500 14500
rect 14600 14400 14700 14500
rect 14800 14400 14900 14500
rect 15000 14400 15100 14500
rect 15200 14400 15300 14500
rect 15400 14400 15500 14500
rect 15600 14400 15700 14500
rect 15800 14400 15900 14500
rect 16000 14400 16100 14500
rect 16200 14400 16300 14500
rect 16400 14400 16500 14500
rect 16600 14400 16700 14500
rect 16800 14400 16900 14500
rect 17000 14400 17100 14500
rect 17200 14400 17300 14500
rect 17400 14400 17500 14500
rect 17600 14400 17700 14500
rect 17800 14400 17900 14500
rect 18000 14400 18100 14500
rect 18200 14400 18300 14500
rect 18400 14400 18500 14500
rect 18600 14400 18700 14500
rect 18800 14400 18900 14500
rect 19000 14400 19100 14500
rect 19200 14400 19300 14500
rect 19400 14400 19500 14500
rect 19600 14400 19700 14500
rect 19800 14400 19900 14500
rect 20000 14400 20100 14500
rect 20200 14400 20300 14500
rect 20400 14400 20500 14500
rect 20600 14400 20700 14500
rect 20800 14400 20900 14500
rect 21000 14400 21100 14500
rect 21200 14400 21300 14500
rect 21400 14400 21500 14500
rect 21600 14400 21700 14500
rect 21800 14400 21900 14500
rect 22000 14400 22100 14500
rect 22200 14400 22300 14500
rect 22400 14400 22500 14500
rect 22600 14400 22700 14500
rect 22800 14400 22900 14500
rect 23000 14400 23100 14500
rect 23200 14400 23300 14500
rect 23400 14400 23500 14500
rect 23600 14400 23700 14500
rect 23800 14400 23900 14500
rect 24000 14400 24100 14500
rect 24200 14400 24300 14500
rect 24400 14400 24500 14500
rect 24600 14400 24700 14500
rect 24800 14400 24900 14500
rect 25000 14400 25100 14500
rect 25200 14400 25300 14500
rect 25400 14400 25500 14500
rect 25600 14400 25700 14500
rect 25800 14400 25900 14500
rect 26000 14400 26100 14500
rect 26200 14400 26300 14500
rect 26400 14400 26500 14500
rect 26600 14400 26700 14500
rect 26800 14400 26900 14500
rect 27000 14400 27100 14500
rect 27200 14400 27300 14500
rect 27400 14400 27500 14500
rect 27600 14400 27700 14500
rect 27800 14400 27900 14500
rect 28000 14400 28100 14500
rect 28200 14400 28300 14500
rect 28400 14400 28500 14500
rect 28600 14400 28700 14500
rect 28800 14400 28900 14500
rect 29000 14400 29100 14500
rect 29200 14400 29300 14500
rect 29400 14400 29500 14500
rect 29600 14400 29700 14500
rect 29800 14400 29900 14500
rect 30000 14400 30100 14500
rect 30200 14400 30300 14500
rect 30400 14400 30500 14500
rect 30600 14400 30700 14500
rect 30800 14400 30900 14500
rect 31000 14400 31100 14500
rect 31200 14400 31300 14500
rect 31400 14400 31500 14500
rect 31600 14400 31700 14500
rect 31800 14400 31900 14500
rect 32000 14400 32100 14500
rect 32200 14400 32300 14500
rect 32400 14400 32500 14500
rect 32600 14400 32700 14500
rect 32800 14400 32900 14500
rect 33000 14400 33100 14500
rect 33200 14400 33316 14500
rect 3200 14300 3300 14400
rect 3200 14100 3300 14200
rect 3200 13900 3300 14000
rect 3200 13700 3300 13800
rect 3200 13500 3300 13600
rect 3200 13300 3300 13400
rect 3200 13100 3300 13200
rect 3200 12900 3300 13000
rect 3200 12700 3300 12800
rect 3200 12500 3300 12600
rect 3200 12300 3300 12400
rect 3200 12100 3300 12200
rect 3200 11900 3300 12000
rect 3200 11700 3300 11800
rect 3200 11500 3300 11600
rect 3200 11300 3300 11400
rect 3200 11100 3300 11200
rect 3200 10900 3300 11000
rect 3200 10700 3300 10800
rect 3200 10500 3300 10600
rect 33200 14300 33300 14400
rect 33200 14100 33300 14200
rect 33200 13900 33300 14000
rect 33200 13700 33300 13800
rect 33200 13500 33300 13600
rect 33200 13300 33300 13400
rect 33200 13100 33300 13200
rect 33200 12900 33300 13000
rect 33200 12700 33300 12800
rect 33200 12500 33300 12600
rect 33200 12300 33300 12400
rect 33200 12100 33300 12200
rect 33200 11900 33300 12000
rect 33200 11700 33300 11800
rect 33200 11500 33300 11600
rect 33200 11300 33300 11400
rect 33200 11100 33300 11200
rect 33200 10900 33300 11000
rect 33200 10700 33300 10800
rect 33200 10500 33300 10600
rect 3184 10400 3300 10500
rect 3400 10400 3500 10500
rect 3600 10400 3700 10500
rect 3800 10400 3900 10500
rect 4000 10400 4100 10500
rect 4200 10400 4300 10500
rect 4400 10400 4500 10500
rect 4600 10400 4700 10500
rect 4800 10400 4900 10500
rect 5000 10400 5100 10500
rect 5200 10400 5300 10500
rect 5400 10400 5500 10500
rect 5600 10400 5700 10500
rect 5800 10400 5900 10500
rect 6000 10400 6100 10500
rect 6200 10400 6300 10500
rect 6400 10400 6500 10500
rect 6600 10400 6700 10500
rect 6800 10400 6900 10500
rect 7000 10400 7100 10500
rect 7200 10400 7300 10500
rect 7400 10400 7500 10500
rect 7600 10400 7700 10500
rect 7800 10400 7900 10500
rect 8000 10400 8100 10500
rect 8200 10400 8300 10500
rect 8400 10400 8500 10500
rect 8600 10400 8700 10500
rect 8800 10400 8900 10500
rect 9000 10400 9100 10500
rect 9200 10400 9300 10500
rect 9400 10400 9500 10500
rect 9600 10400 9700 10500
rect 9800 10400 9900 10500
rect 10000 10400 10100 10500
rect 10200 10400 10300 10500
rect 10400 10400 10500 10500
rect 10600 10400 10700 10500
rect 10800 10400 10900 10500
rect 11000 10400 11100 10500
rect 11200 10400 11300 10500
rect 11400 10400 11500 10500
rect 11600 10400 11700 10500
rect 11800 10400 11900 10500
rect 12000 10400 12100 10500
rect 12200 10400 12300 10500
rect 12400 10400 12500 10500
rect 12600 10400 12700 10500
rect 12800 10400 12900 10500
rect 13000 10400 13100 10500
rect 13200 10400 13300 10500
rect 13400 10400 13500 10500
rect 13600 10400 13700 10500
rect 13800 10400 13900 10500
rect 14000 10400 14100 10500
rect 14200 10400 14300 10500
rect 14400 10400 14500 10500
rect 14600 10400 14700 10500
rect 14800 10400 14900 10500
rect 15000 10400 15100 10500
rect 15200 10400 15300 10500
rect 15400 10400 15500 10500
rect 15600 10400 15700 10500
rect 15800 10400 15900 10500
rect 16000 10400 16100 10500
rect 16200 10400 16300 10500
rect 16400 10400 16500 10500
rect 16600 10400 16700 10500
rect 16800 10400 16900 10500
rect 17000 10400 17100 10500
rect 17200 10400 17300 10500
rect 17400 10400 17500 10500
rect 17600 10400 17700 10500
rect 17800 10400 17900 10500
rect 18000 10400 18100 10500
rect 18200 10400 18300 10500
rect 18400 10400 18500 10500
rect 18600 10400 18700 10500
rect 18800 10400 18900 10500
rect 19000 10400 19100 10500
rect 19200 10400 19300 10500
rect 19400 10400 19500 10500
rect 19600 10400 19700 10500
rect 19800 10400 19900 10500
rect 20000 10400 20100 10500
rect 20200 10400 20300 10500
rect 20400 10400 20500 10500
rect 20600 10400 20700 10500
rect 20800 10400 20900 10500
rect 21000 10400 21100 10500
rect 21200 10400 21300 10500
rect 21400 10400 21500 10500
rect 21600 10400 21700 10500
rect 21800 10400 21900 10500
rect 22000 10400 22100 10500
rect 22200 10400 22300 10500
rect 22400 10400 22500 10500
rect 22600 10400 22700 10500
rect 22800 10400 22900 10500
rect 23000 10400 23100 10500
rect 23200 10400 23300 10500
rect 23400 10400 23500 10500
rect 23600 10400 23700 10500
rect 23800 10400 23900 10500
rect 24000 10400 24100 10500
rect 24200 10400 24300 10500
rect 24400 10400 24500 10500
rect 24600 10400 24700 10500
rect 24800 10400 24900 10500
rect 25000 10400 25100 10500
rect 25200 10400 25300 10500
rect 25400 10400 25500 10500
rect 25600 10400 25700 10500
rect 25800 10400 25900 10500
rect 26000 10400 26100 10500
rect 26200 10400 26300 10500
rect 26400 10400 26500 10500
rect 26600 10400 26700 10500
rect 26800 10400 26900 10500
rect 27000 10400 27100 10500
rect 27200 10400 27300 10500
rect 27400 10400 27500 10500
rect 27600 10400 27700 10500
rect 27800 10400 27900 10500
rect 28000 10400 28100 10500
rect 28200 10400 28300 10500
rect 28400 10400 28500 10500
rect 28600 10400 28700 10500
rect 28800 10400 28900 10500
rect 29000 10400 29100 10500
rect 29200 10400 29300 10500
rect 29400 10400 29500 10500
rect 29600 10400 29700 10500
rect 29800 10400 29900 10500
rect 30000 10400 30100 10500
rect 30200 10400 30300 10500
rect 30400 10400 30500 10500
rect 30600 10400 30700 10500
rect 30800 10400 30900 10500
rect 31000 10400 31100 10500
rect 31200 10400 31300 10500
rect 31400 10400 31500 10500
rect 31600 10400 31700 10500
rect 31800 10400 31900 10500
rect 32000 10400 32100 10500
rect 32200 10400 32300 10500
rect 32400 10400 32500 10500
rect 32600 10400 32700 10500
rect 32800 10400 32900 10500
rect 33000 10400 33100 10500
rect 33200 10400 33316 10500
rect 184 10000 300 10100
rect 400 10000 500 10100
rect 600 10000 700 10100
rect 800 10000 900 10100
rect 1000 10000 1100 10100
rect 1200 10000 1300 10100
rect 1400 10000 1500 10100
rect 1600 10000 1700 10100
rect 1800 10000 1900 10100
rect 2000 10000 2100 10100
rect 2200 10000 2300 10100
rect 2400 10000 2500 10100
rect 2600 10000 2700 10100
rect 2800 10000 2900 10100
rect 3000 10000 3100 10100
rect 3200 10000 3300 10100
rect 3400 10000 3500 10100
rect 3600 10000 3700 10100
rect 3800 10000 3900 10100
rect 4000 10000 4100 10100
rect 4200 10000 4300 10100
rect 4400 10000 4500 10100
rect 4600 10000 4700 10100
rect 4800 10000 4900 10100
rect 5000 10000 5100 10100
rect 5200 10000 5300 10100
rect 5400 10000 5500 10100
rect 5600 10000 5700 10100
rect 5800 10000 5900 10100
rect 6000 10000 6100 10100
rect 6200 10000 6300 10100
rect 6400 10000 6500 10100
rect 6600 10000 6700 10100
rect 6800 10000 6900 10100
rect 7000 10000 7100 10100
rect 7200 10000 7300 10100
rect 7400 10000 7500 10100
rect 7600 10000 7700 10100
rect 7800 10000 7900 10100
rect 8000 10000 8100 10100
rect 8200 10000 8300 10100
rect 8400 10000 8500 10100
rect 8600 10000 8700 10100
rect 8800 10000 8900 10100
rect 9000 10000 9100 10100
rect 9200 10000 9300 10100
rect 9400 10000 9500 10100
rect 9600 10000 9700 10100
rect 9800 10000 9900 10100
rect 10000 10000 10100 10100
rect 10200 10000 10300 10100
rect 10400 10000 10500 10100
rect 10600 10000 10700 10100
rect 10800 10000 10900 10100
rect 11000 10000 11100 10100
rect 11200 10000 11300 10100
rect 11400 10000 11500 10100
rect 11600 10000 11700 10100
rect 11800 10000 11900 10100
rect 12000 10000 12100 10100
rect 12200 10000 12300 10100
rect 12400 10000 12500 10100
rect 12600 10000 12700 10100
rect 12800 10000 12900 10100
rect 13000 10000 13100 10100
rect 13200 10000 13300 10100
rect 13400 10000 13500 10100
rect 13600 10000 13700 10100
rect 13800 10000 13900 10100
rect 14000 10000 14100 10100
rect 14200 10000 14300 10100
rect 14400 10000 14500 10100
rect 14600 10000 14700 10100
rect 14800 10000 14900 10100
rect 15000 10000 15100 10100
rect 15200 10000 15300 10100
rect 15400 10000 15500 10100
rect 15600 10000 15700 10100
rect 15800 10000 15900 10100
rect 16000 10000 16100 10100
rect 16200 10000 16300 10100
rect 16400 10000 16500 10100
rect 16600 10000 16700 10100
rect 16800 10000 16900 10100
rect 17000 10000 17100 10100
rect 17200 10000 17300 10100
rect 17400 10000 17500 10100
rect 17600 10000 17700 10100
rect 17800 10000 17900 10100
rect 18000 10000 18100 10100
rect 18200 10000 18300 10100
rect 18400 10000 18500 10100
rect 18600 10000 18700 10100
rect 18800 10000 18900 10100
rect 19000 10000 19100 10100
rect 19200 10000 19300 10100
rect 19400 10000 19500 10100
rect 19600 10000 19700 10100
rect 19800 10000 19900 10100
rect 20000 10000 20100 10100
rect 20200 10000 20300 10100
rect 20400 10000 20500 10100
rect 20600 10000 20700 10100
rect 20800 10000 20900 10100
rect 21000 10000 21100 10100
rect 21200 10000 21300 10100
rect 21400 10000 21500 10100
rect 21600 10000 21700 10100
rect 21800 10000 21900 10100
rect 22000 10000 22100 10100
rect 22200 10000 22300 10100
rect 22400 10000 22500 10100
rect 22600 10000 22700 10100
rect 22800 10000 22900 10100
rect 23000 10000 23100 10100
rect 23200 10000 23300 10100
rect 23400 10000 23500 10100
rect 23600 10000 23700 10100
rect 23800 10000 23900 10100
rect 24000 10000 24100 10100
rect 24200 10000 24300 10100
rect 24400 10000 24500 10100
rect 24600 10000 24700 10100
rect 24800 10000 24900 10100
rect 25000 10000 25100 10100
rect 25200 10000 25300 10100
rect 25400 10000 25500 10100
rect 25600 10000 25700 10100
rect 25800 10000 25900 10100
rect 26000 10000 26100 10100
rect 26200 10000 26300 10100
rect 26400 10000 26500 10100
rect 26600 10000 26700 10100
rect 26800 10000 26900 10100
rect 27000 10000 27100 10100
rect 27200 10000 27300 10100
rect 27400 10000 27500 10100
rect 27600 10000 27700 10100
rect 27800 10000 27900 10100
rect 28000 10000 28100 10100
rect 28200 10000 28300 10100
rect 28400 10000 28500 10100
rect 28600 10000 28700 10100
rect 28800 10000 28900 10100
rect 29000 10000 29100 10100
rect 29200 10000 29300 10100
rect 29400 10000 29500 10100
rect 29600 10000 29700 10100
rect 29800 10000 29900 10100
rect 30000 10000 30100 10100
rect 30200 10000 30300 10100
rect 30400 10000 30500 10100
rect 30600 10000 30700 10100
rect 30800 10000 30900 10100
rect 31000 10000 31100 10100
rect 31200 10000 31300 10100
rect 31400 10000 31500 10100
rect 31600 10000 31700 10100
rect 31800 10000 31900 10100
rect 32000 10000 32100 10100
rect 32200 10000 32300 10100
rect 32400 10000 32500 10100
rect 32600 10000 32700 10100
rect 32800 10000 32900 10100
rect 33000 10000 33100 10100
rect 33200 10000 33300 10100
rect 33400 10000 33500 10100
rect 33600 10000 33700 10100
rect 33800 10000 33900 10100
rect 34000 10000 34100 10100
rect 34200 10000 34300 10100
rect 34400 10000 34500 10100
rect 34600 10000 34700 10100
rect 34800 10000 34900 10100
rect 35000 10000 35100 10100
rect 35200 10000 35300 10100
rect 35400 10000 35500 10100
rect 35600 10000 35700 10100
rect 35800 10000 35900 10100
rect 36000 10000 36116 10100
rect 200 9900 300 10000
rect 200 9700 300 9800
rect 200 9500 300 9600
rect 200 9300 300 9400
rect 200 9100 300 9200
rect 200 8900 300 9000
rect 200 8700 300 8800
rect 200 8500 300 8600
rect 200 8300 300 8400
rect 200 8100 300 8200
rect 200 7900 300 8000
rect 200 7700 300 7800
rect 200 7500 300 7600
rect 200 7300 300 7400
rect 200 7100 300 7200
rect 200 6900 300 7000
rect 200 6700 300 6800
rect 200 6500 300 6600
rect 200 6300 300 6400
rect 200 6100 300 6200
rect 36000 9900 36100 10000
rect 36000 9700 36100 9800
rect 36000 9500 36100 9600
rect 36000 9300 36100 9400
rect 36000 9100 36100 9200
rect 36000 8900 36100 9000
rect 36000 8700 36100 8800
rect 36000 8500 36100 8600
rect 36000 8300 36100 8400
rect 36000 8100 36100 8200
rect 36000 7900 36100 8000
rect 36000 7700 36100 7800
rect 36000 7500 36100 7600
rect 36000 7300 36100 7400
rect 36000 7100 36100 7200
rect 36000 6900 36100 7000
rect 36000 6700 36100 6800
rect 36000 6500 36100 6600
rect 36000 6300 36100 6400
rect 36000 6100 36100 6200
rect 184 6000 300 6100
rect 400 6000 500 6100
rect 600 6000 700 6100
rect 800 6000 900 6100
rect 1000 6000 1100 6100
rect 1200 6000 1300 6100
rect 1400 6000 1500 6100
rect 1600 6000 1700 6100
rect 1800 6000 1900 6100
rect 2000 6000 2100 6100
rect 2200 6000 2300 6100
rect 2400 6000 2500 6100
rect 2600 6000 2700 6100
rect 2800 6000 2900 6100
rect 3000 6000 3100 6100
rect 3200 6000 3300 6100
rect 3400 6000 3500 6100
rect 3600 6000 3700 6100
rect 3800 6000 3900 6100
rect 4000 6000 4100 6100
rect 4200 6000 4300 6100
rect 4400 6000 4500 6100
rect 4600 6000 4700 6100
rect 4800 6000 4900 6100
rect 5000 6000 5100 6100
rect 5200 6000 5300 6100
rect 5400 6000 5500 6100
rect 5600 6000 5700 6100
rect 5800 6000 5900 6100
rect 6000 6000 6100 6100
rect 6200 6000 6300 6100
rect 6400 6000 6500 6100
rect 6600 6000 6700 6100
rect 6800 6000 6900 6100
rect 7000 6000 7100 6100
rect 7200 6000 7300 6100
rect 7400 6000 7500 6100
rect 7600 6000 7700 6100
rect 7800 6000 7900 6100
rect 8000 6000 8100 6100
rect 8200 6000 8300 6100
rect 8400 6000 8500 6100
rect 8600 6000 8700 6100
rect 8800 6000 8900 6100
rect 9000 6000 9100 6100
rect 9200 6000 9300 6100
rect 9400 6000 9500 6100
rect 9600 6000 9700 6100
rect 9800 6000 9900 6100
rect 10000 6000 10100 6100
rect 10200 6000 10300 6100
rect 10400 6000 10500 6100
rect 10600 6000 10700 6100
rect 10800 6000 10900 6100
rect 11000 6000 11100 6100
rect 11200 6000 11300 6100
rect 11400 6000 11500 6100
rect 11600 6000 11700 6100
rect 11800 6000 11900 6100
rect 12000 6000 12100 6100
rect 12200 6000 12300 6100
rect 12400 6000 12500 6100
rect 12600 6000 12700 6100
rect 12800 6000 12900 6100
rect 13000 6000 13100 6100
rect 13200 6000 13300 6100
rect 13400 6000 13500 6100
rect 13600 6000 13700 6100
rect 13800 6000 13900 6100
rect 14000 6000 14100 6100
rect 14200 6000 14300 6100
rect 14400 6000 14500 6100
rect 14600 6000 14700 6100
rect 14800 6000 14900 6100
rect 15000 6000 15100 6100
rect 15200 6000 15300 6100
rect 15400 6000 15500 6100
rect 15600 6000 15700 6100
rect 15800 6000 15900 6100
rect 16000 6000 16100 6100
rect 16200 6000 16300 6100
rect 16400 6000 16500 6100
rect 16600 6000 16700 6100
rect 16800 6000 16900 6100
rect 17000 6000 17100 6100
rect 17200 6000 17300 6100
rect 17400 6000 17500 6100
rect 17600 6000 17700 6100
rect 17800 6000 17900 6100
rect 18000 6000 18100 6100
rect 18200 6000 18300 6100
rect 18400 6000 18500 6100
rect 18600 6000 18700 6100
rect 18800 6000 18900 6100
rect 19000 6000 19100 6100
rect 19200 6000 19300 6100
rect 19400 6000 19500 6100
rect 19600 6000 19700 6100
rect 19800 6000 19900 6100
rect 20000 6000 20100 6100
rect 20200 6000 20300 6100
rect 20400 6000 20500 6100
rect 20600 6000 20700 6100
rect 20800 6000 20900 6100
rect 21000 6000 21100 6100
rect 21200 6000 21300 6100
rect 21400 6000 21500 6100
rect 21600 6000 21700 6100
rect 21800 6000 21900 6100
rect 22000 6000 22100 6100
rect 22200 6000 22300 6100
rect 22400 6000 22500 6100
rect 22600 6000 22700 6100
rect 22800 6000 22900 6100
rect 23000 6000 23100 6100
rect 23200 6000 23300 6100
rect 23400 6000 23500 6100
rect 23600 6000 23700 6100
rect 23800 6000 23900 6100
rect 24000 6000 24100 6100
rect 24200 6000 24300 6100
rect 24400 6000 24500 6100
rect 24600 6000 24700 6100
rect 24800 6000 24900 6100
rect 25000 6000 25100 6100
rect 25200 6000 25300 6100
rect 25400 6000 25500 6100
rect 25600 6000 25700 6100
rect 25800 6000 25900 6100
rect 26000 6000 26100 6100
rect 26200 6000 26300 6100
rect 26400 6000 26500 6100
rect 26600 6000 26700 6100
rect 26800 6000 26900 6100
rect 27000 6000 27100 6100
rect 27200 6000 27300 6100
rect 27400 6000 27500 6100
rect 27600 6000 27700 6100
rect 27800 6000 27900 6100
rect 28000 6000 28100 6100
rect 28200 6000 28300 6100
rect 28400 6000 28500 6100
rect 28600 6000 28700 6100
rect 28800 6000 28900 6100
rect 29000 6000 29100 6100
rect 29200 6000 29300 6100
rect 29400 6000 29500 6100
rect 29600 6000 29700 6100
rect 29800 6000 29900 6100
rect 30000 6000 30100 6100
rect 30200 6000 30300 6100
rect 30400 6000 30500 6100
rect 30600 6000 30700 6100
rect 30800 6000 30900 6100
rect 31000 6000 31100 6100
rect 31200 6000 31300 6100
rect 31400 6000 31500 6100
rect 31600 6000 31700 6100
rect 31800 6000 31900 6100
rect 32000 6000 32100 6100
rect 32200 6000 32300 6100
rect 32400 6000 32500 6100
rect 32600 6000 32700 6100
rect 32800 6000 32900 6100
rect 33000 6000 33100 6100
rect 33200 6000 33300 6100
rect 33400 6000 33500 6100
rect 33600 6000 33700 6100
rect 33800 6000 33900 6100
rect 34000 6000 34100 6100
rect 34200 6000 34300 6100
rect 34400 6000 34500 6100
rect 34600 6000 34700 6100
rect 34800 6000 34900 6100
rect 35000 6000 35100 6100
rect 35200 6000 35300 6100
rect 35400 6000 35500 6100
rect 35600 6000 35700 6100
rect 35800 6000 35900 6100
rect 36000 6000 36116 6100
<< labels >>
flabel locali 32246 10400 32636 10500 1 FreeSans 1600 0 0 0 gnd
flabel locali 32253 10000 32643 10100 1 FreeSans 1600 0 0 0 gnd
<< end >>
