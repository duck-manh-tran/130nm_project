* SPICE3 file created from vco_w6_r100.ext - technology: sky130A
*input_sig enb vdd gnd v_ctr
.subckt vco_w6_r100 p[0] p[1] p[3] p[5] p[7] p[9] p[10] p[8] p[6] p[4] p[2] input_analog enb vccd2 vssd2 
R0 ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__res_generic_po w=2 l=4.15
R1 ring_osc_w6_0/v_ctr input_analog sky130_fd_pr__res_generic_po w=2 l=4.15
X0 vccd2 p[8] p[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X1 p[10] p[8] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X2 vccd2 ring_osc_w6_0/pn[9] ring_osc_w6_0/pn[10] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X3 ring_osc_w6_0/pn[10] ring_osc_w6_0/pn[9] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X4 ring_osc_w6_0/pn[10] p[10] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X5 p[10] ring_osc_w6_0/pn[10] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X6 ring_osc_w6_0/v_ctr p[8] p[10] ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X7 p[10] p[8] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X8 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[9] ring_osc_w6_0/pn[10] ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X9 ring_osc_w6_0/pn[10] ring_osc_w6_0/pn[9] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_10/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X10 ring_osc_w6_0/pn[10] p[10] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X11 p[10] ring_osc_w6_0/pn[10] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X12 vccd2 p[10] p[9] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X13 p[9] p[10] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X14 vccd2 ring_osc_w6_0/pn[10] ring_osc_w6_0/pn[0] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X15 ring_osc_w6_0/pn[0] ring_osc_w6_0/pn[10] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X16 ring_osc_w6_0/pn[0] p[9] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X17 p[9] ring_osc_w6_0/pn[0] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X18 ring_osc_w6_0/v_ctr p[10] p[9] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X19 p[9] p[10] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X20 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[10] ring_osc_w6_0/pn[0] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X21 ring_osc_w6_0/pn[0] ring_osc_w6_0/pn[10] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X22 ring_osc_w6_0/pn[0] p[9] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X23 p[9] ring_osc_w6_0/pn[0] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X24 vccd2 p[9] p[7] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X25 p[7] p[9] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X26 vccd2 ring_osc_w6_0/pn[0] ring_osc_w6_0/pn[1] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X27 ring_osc_w6_0/pn[1] ring_osc_w6_0/pn[0] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X28 ring_osc_w6_0/pn[1] p[7] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X29 p[7] ring_osc_w6_0/pn[1] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X30 ring_osc_w6_0/v_ctr p[9] p[7] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X31 p[7] p[9] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X32 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[0] ring_osc_w6_0/pn[1] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X33 ring_osc_w6_0/pn[1] ring_osc_w6_0/pn[0] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X34 ring_osc_w6_0/pn[1] p[7] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X35 p[7] ring_osc_w6_0/pn[1] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X36 vccd2 p[7] p[5] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X37 p[5] p[7] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X38 vccd2 ring_osc_w6_0/pn[1] ring_osc_w6_0/pn[2] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X39 ring_osc_w6_0/pn[2] ring_osc_w6_0/pn[1] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X40 ring_osc_w6_0/pn[2] p[5] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X41 p[5] ring_osc_w6_0/pn[2] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X42 ring_osc_w6_0/v_ctr p[7] p[5] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X43 p[5] p[7] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X44 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[1] ring_osc_w6_0/pn[2] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X45 ring_osc_w6_0/pn[2] ring_osc_w6_0/pn[1] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X46 ring_osc_w6_0/pn[2] p[5] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X47 p[5] ring_osc_w6_0/pn[2] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
R2 ring_osc_w6_0/sky130_fd_sc_hd__einvp_1_0/A vccd2 sky130_fd_pr__res_generic_po w=480000u l=45000u
R3 vssd2 ring_osc_w6_0/sky130_fd_sc_hd__conb_1_0/LO sky130_fd_pr__res_generic_po w=480000u l=45000u
X48 vccd2 p[5] p[3] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X49 p[3] p[5] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X50 vccd2 ring_osc_w6_0/pn[2] ring_osc_w6_0/pn[3] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X51 ring_osc_w6_0/pn[3] ring_osc_w6_0/pn[2] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X52 ring_osc_w6_0/pn[3] p[3] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X53 p[3] ring_osc_w6_0/pn[3] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X54 ring_osc_w6_0/v_ctr p[5] p[3] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X55 p[3] p[5] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X56 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[2] ring_osc_w6_0/pn[3] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X57 ring_osc_w6_0/pn[3] ring_osc_w6_0/pn[2] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X58 ring_osc_w6_0/pn[3] p[3] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X59 p[3] ring_osc_w6_0/pn[3] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X60 vccd2 p[3] p[1] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X61 p[1] p[3] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X62 vccd2 ring_osc_w6_0/pn[3] ring_osc_w6_0/pn[4] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X63 ring_osc_w6_0/pn[4] ring_osc_w6_0/pn[3] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X64 ring_osc_w6_0/pn[4] p[1] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X65 p[1] ring_osc_w6_0/pn[4] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X66 ring_osc_w6_0/v_ctr p[3] p[1] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X67 p[1] p[3] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X68 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[3] ring_osc_w6_0/pn[4] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X69 ring_osc_w6_0/pn[4] ring_osc_w6_0/pn[3] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X70 ring_osc_w6_0/pn[4] p[1] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X71 p[1] ring_osc_w6_0/pn[4] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X72 vccd2 p[1] p[0] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X73 p[0] p[1] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X74 vccd2 ring_osc_w6_0/pn[4] ring_osc_w6_0/pn[5] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X75 ring_osc_w6_0/pn[5] ring_osc_w6_0/pn[4] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X76 ring_osc_w6_0/pn[5] p[0] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X77 p[0] ring_osc_w6_0/pn[5] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X78 ring_osc_w6_0/v_ctr p[1] p[0] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X79 p[0] p[1] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X80 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[4] ring_osc_w6_0/pn[5] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X81 ring_osc_w6_0/pn[5] ring_osc_w6_0/pn[4] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X82 ring_osc_w6_0/pn[5] p[0] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X83 p[0] ring_osc_w6_0/pn[5] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X84 vccd2 p[2] p[4] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X85 p[4] p[2] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X86 vccd2 ring_osc_w6_0/pn[6] ring_osc_w6_0/pn[7] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X87 ring_osc_w6_0/pn[7] ring_osc_w6_0/pn[6] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X88 ring_osc_w6_0/pn[7] p[4] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X89 p[4] ring_osc_w6_0/pn[7] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X90 ring_osc_w6_0/v_ctr p[2] p[4] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X91 p[4] p[2] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X92 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[6] ring_osc_w6_0/pn[7] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X93 ring_osc_w6_0/pn[7] ring_osc_w6_0/pn[6] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X94 ring_osc_w6_0/pn[7] p[4] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X95 p[4] ring_osc_w6_0/pn[7] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X96 vccd2 p[0] p[2] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X97 p[2] p[0] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X98 vccd2 ring_osc_w6_0/pn[5] ring_osc_w6_0/pn[6] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X99 ring_osc_w6_0/pn[6] ring_osc_w6_0/pn[5] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X100 ring_osc_w6_0/pn[6] p[2] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X101 p[2] ring_osc_w6_0/pn[6] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X102 ring_osc_w6_0/v_ctr p[0] p[2] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X103 p[2] p[0] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X104 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[5] ring_osc_w6_0/pn[6] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X105 ring_osc_w6_0/pn[6] ring_osc_w6_0/pn[5] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X106 ring_osc_w6_0/pn[6] p[2] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X107 p[2] ring_osc_w6_0/pn[6] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X108 vccd2 p[4] p[6] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X109 p[6] p[4] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X110 vccd2 ring_osc_w6_0/pn[7] ring_osc_w6_0/pn[8] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X111 ring_osc_w6_0/pn[8] ring_osc_w6_0/pn[7] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X112 ring_osc_w6_0/pn[8] p[6] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X113 p[6] ring_osc_w6_0/pn[8] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X114 ring_osc_w6_0/v_ctr p[4] p[6] ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X115 p[6] p[4] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X116 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[7] ring_osc_w6_0/pn[8] ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X117 ring_osc_w6_0/pn[8] ring_osc_w6_0/pn[7] ring_osc_w6_0/v_ctr ring_osc_w6_0/inv_8/vssd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X118 ring_osc_w6_0/pn[8] p[6] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X119 p[6] ring_osc_w6_0/pn[8] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X120 vccd2 p[6] p[8] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X121 p[8] p[6] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X122 vccd2 ring_osc_w6_0/pn[8] ring_osc_w6_0/pn[9] vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X123 ring_osc_w6_0/pn[9] ring_osc_w6_0/pn[8] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X124 ring_osc_w6_0/pn[9] p[8] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X125 p[8] ring_osc_w6_0/pn[9] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X126 ring_osc_w6_0/v_ctr p[6] p[8] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X127 p[8] p[6] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X128 ring_osc_w6_0/v_ctr ring_osc_w6_0/pn[8] ring_osc_w6_0/pn[9] vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X129 ring_osc_w6_0/pn[9] ring_osc_w6_0/pn[8] ring_osc_w6_0/v_ctr vssd2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X130 ring_osc_w6_0/pn[9] p[8] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X131 p[8] ring_osc_w6_0/pn[9] vccd2 vccd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5 l=1.9
X132 a_1627_12582# li_1496_12384# vccd2 vccd2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1 l=150000u
X133 p[0] ring_osc_w6_0/sky130_fd_sc_hd__einvp_1_0/A a_1627_12258# ring_osc_w6_0/sky130_fd_sc_hd__conb_1_0/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=-0p ps=0u w=650000u l=150000u
X134 vccd2 enb li_1496_12384# vccd2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X135 p[0] ring_osc_w6_0/sky130_fd_sc_hd__einvp_1_0/A a_1627_12582# vccd2 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1 l=150000u
X136 a_1627_12258# enb vssd2 ring_osc_w6_0/sky130_fd_sc_hd__conb_1_0/VNB sky130_fd_pr__nfet_01v8 ad=-0p pd=0u as=0p ps=0u w=650000u l=150000u
X137 vssd2 enb li_1496_12384# ring_osc_w6_0/sky130_fd_sc_hd__conb_1_0/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 ring_osc_w6_0/pn[10] p[10] 3.59fF
C1 p[2] vccd2 2.80fF
C2 vccd2 p[5] 2.64fF
C3 p[2] ring_osc_w6_0/pn[6] 2.82fF
C4 p[3] ring_osc_w6_0/pn[3] 2.51fF
C5 ring_osc_w6_0/pn[5] ring_osc_w6_0/v_ctr 2.54fF
C6 ring_osc_w6_0/pn[1] p[7] 2.52fF
C7 ring_osc_w6_0/pn[2] p[5] 2.73fF
C8 vccd2 p[0] 3.44fF
C9 p[8] ring_osc_w6_0/pn[9] 2.78fF
C10 p[9] ring_osc_w6_0/pn[0] 2.91fF
C11 ring_osc_w6_0/pn[4] vccd2 2.26fF
C12 ring_osc_w6_0/pn[10] ring_osc_w6_0/v_ctr 2.65fF
C13 ring_osc_w6_0/pn[5] p[0] 3.56fF
C14 vccd2 p[6] 2.82fF
C15 ring_osc_w6_0/pn[7] p[4] 2.73fF
C16 vccd2 ring_osc_w6_0/pn[8] 2.09fF
C17 p[6] ring_osc_w6_0/pn[8] 2.73fF
C18 vccd2 p[7] 3.66fF
C19 vccd2 p[9] 2.94fF
C20 ring_osc_w6_0/pn[4] p[1] 2.28fF
C21 vccd2 p[1] 2.36fF
C22 p[8] vccd2 2.35fF
C23 vccd2 ring_osc_w6_0/pn[10] 2.95fF
C24 p[3] vccd2 3.07fF
C25 vccd2 p[4] 3.18fF
C26 vccd2 ring_osc_w6_0/v_ctr 6.18fF
C27 vccd2 ring_osc_w6_0/sky130_fd_sc_hd__conb_1_0/VNB 363.00fF
.ends
