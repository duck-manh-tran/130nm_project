* Subcircuit       : ring_osc
* Library          : ADC_130nm
* Generate for     : NGSPICE (ngbehavior=hs)
********************************************************************************
.subckt ring_osc vdd vss 
+ p[0] p[1] p[2] p[3] p[4] p[5] p[6] p[7] p[8] p[9] p[10]
+ Ln12=0.36 Wn12=1 Fn12=1 Lp12=0.36 Wp12=1 Fp12=1
+ Ln34=0.36 Wn34=1 Fn34=1 Lp34=0.36 Wp34=1 Fp34=1

*phase0_inv0(out -> p[0])
Xc1 p[10] p_n[10] p[0] p_n[0] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34


*phase1_inv1(out -> p[1])
Xc2 p[0] p_n[0] p[1] p_n[1] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv2(out -> p[2])
Xc3 p[1] p_n[1] p[2] p_n[2] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv3(out -> p[3])
Xc4 p[2] p_n[2] p[3] p_n[3] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv4(out -> p[4])
Xc5 p[3] p_n[3] p[4] p_n[4] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv5(out -> p[5])
Xc6 p[4] p_n[4] p[5] p_n[5] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv6(out -> p[6])
Xc7 p[5] p_n[5] p[6] p_n[6] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv7(out -> p[7])
Xc8 p[6] p_n[6] p[7] p_n[7] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv8(out -> p[8])
Xc9 p[7] p_n[7] p[8] p_n[8] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv9(out -> p[9])
Xc10 p[8] p_n[8] p[9] p_n[9] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34



*phase1_inv10(out -> p[10])
Xc11 p[9] p_n[9] p[10] p_n[10] vdd vss crs_cpl_inv
+ Ln_12=Ln12 Wn_12=Wn12 Fn_12=Fn12 Lp_12=Lp12 Wp_12=Wp12 Fp_12=Fp12
+ Ln_34=Ln34 Wn_34=Wn34 Fn_34=Fn34 Lp_34=Lp34 Wp_34=Wp34 Fp_34=Fp34


.ends ring_osc


*note:
* .subckt crs_cpl_inv inp inn outp outn vdd vss
* + Ln_12=0.36 Wn_12=1 Fn_12=1 Lp_12=0.36 Wp_12=1 Fp_12=1
* + Ln_34=0.36 Wn_34=1 Fn_34=1 Lp_34=0.36 Wp_34=1 Fp_34=1

