magic
tech sky130A
timestamp 1637143825
<< nwell >>
rect 0 0 700 1000
<< pmos >>
rect 145 100 335 900
rect 365 100 555 900
<< pdiff >>
rect 115 887 145 900
rect 115 869 121 887
rect 139 869 145 887
rect 115 851 145 869
rect 115 833 121 851
rect 139 833 145 851
rect 115 815 145 833
rect 115 797 121 815
rect 139 797 145 815
rect 115 779 145 797
rect 115 761 121 779
rect 139 761 145 779
rect 115 743 145 761
rect 115 725 121 743
rect 139 725 145 743
rect 115 707 145 725
rect 115 689 121 707
rect 139 689 145 707
rect 115 671 145 689
rect 115 653 121 671
rect 139 653 145 671
rect 115 635 145 653
rect 115 617 121 635
rect 139 617 145 635
rect 115 599 145 617
rect 115 581 121 599
rect 139 581 145 599
rect 115 563 145 581
rect 115 545 121 563
rect 139 545 145 563
rect 115 527 145 545
rect 115 509 121 527
rect 139 509 145 527
rect 115 491 145 509
rect 115 473 121 491
rect 139 473 145 491
rect 115 455 145 473
rect 115 437 121 455
rect 139 437 145 455
rect 115 419 145 437
rect 115 401 121 419
rect 139 401 145 419
rect 115 383 145 401
rect 115 365 121 383
rect 139 365 145 383
rect 115 347 145 365
rect 115 329 121 347
rect 139 329 145 347
rect 115 311 145 329
rect 115 293 121 311
rect 139 293 145 311
rect 115 275 145 293
rect 115 257 121 275
rect 139 257 145 275
rect 115 239 145 257
rect 115 221 121 239
rect 139 221 145 239
rect 115 203 145 221
rect 115 185 121 203
rect 139 185 145 203
rect 115 167 145 185
rect 115 149 121 167
rect 139 149 145 167
rect 115 131 145 149
rect 115 113 121 131
rect 139 113 145 131
rect 115 100 145 113
rect 335 887 365 900
rect 335 869 341 887
rect 359 869 365 887
rect 335 851 365 869
rect 335 833 341 851
rect 359 833 365 851
rect 335 815 365 833
rect 335 797 341 815
rect 359 797 365 815
rect 335 779 365 797
rect 335 761 341 779
rect 359 761 365 779
rect 335 743 365 761
rect 335 725 341 743
rect 359 725 365 743
rect 335 707 365 725
rect 335 689 341 707
rect 359 689 365 707
rect 335 671 365 689
rect 335 653 341 671
rect 359 653 365 671
rect 335 635 365 653
rect 335 617 341 635
rect 359 617 365 635
rect 335 599 365 617
rect 335 581 341 599
rect 359 581 365 599
rect 335 563 365 581
rect 335 545 341 563
rect 359 545 365 563
rect 335 527 365 545
rect 335 509 341 527
rect 359 509 365 527
rect 335 491 365 509
rect 335 473 341 491
rect 359 473 365 491
rect 335 455 365 473
rect 335 437 341 455
rect 359 437 365 455
rect 335 419 365 437
rect 335 401 341 419
rect 359 401 365 419
rect 335 383 365 401
rect 335 365 341 383
rect 359 365 365 383
rect 335 347 365 365
rect 335 329 341 347
rect 359 329 365 347
rect 335 311 365 329
rect 335 293 341 311
rect 359 293 365 311
rect 335 275 365 293
rect 335 257 341 275
rect 359 257 365 275
rect 335 239 365 257
rect 335 221 341 239
rect 359 221 365 239
rect 335 203 365 221
rect 335 185 341 203
rect 359 185 365 203
rect 335 167 365 185
rect 335 149 341 167
rect 359 149 365 167
rect 335 131 365 149
rect 335 113 341 131
rect 359 113 365 131
rect 335 100 365 113
rect 555 887 585 900
rect 555 869 561 887
rect 579 869 585 887
rect 555 851 585 869
rect 555 833 561 851
rect 579 833 585 851
rect 555 815 585 833
rect 555 797 561 815
rect 579 797 585 815
rect 555 779 585 797
rect 555 761 561 779
rect 579 761 585 779
rect 555 743 585 761
rect 555 725 561 743
rect 579 725 585 743
rect 555 707 585 725
rect 555 689 561 707
rect 579 689 585 707
rect 555 671 585 689
rect 555 653 561 671
rect 579 653 585 671
rect 555 635 585 653
rect 555 617 561 635
rect 579 617 585 635
rect 555 599 585 617
rect 555 581 561 599
rect 579 581 585 599
rect 555 563 585 581
rect 555 545 561 563
rect 579 545 585 563
rect 555 527 585 545
rect 555 509 561 527
rect 579 509 585 527
rect 555 491 585 509
rect 555 473 561 491
rect 579 473 585 491
rect 555 455 585 473
rect 555 437 561 455
rect 579 437 585 455
rect 555 419 585 437
rect 555 401 561 419
rect 579 401 585 419
rect 555 383 585 401
rect 555 365 561 383
rect 579 365 585 383
rect 555 347 585 365
rect 555 329 561 347
rect 579 329 585 347
rect 555 311 585 329
rect 555 293 561 311
rect 579 293 585 311
rect 555 275 585 293
rect 555 257 561 275
rect 579 257 585 275
rect 555 239 585 257
rect 555 221 561 239
rect 579 221 585 239
rect 555 203 585 221
rect 555 185 561 203
rect 579 185 585 203
rect 555 167 585 185
rect 555 149 561 167
rect 579 149 585 167
rect 555 131 585 149
rect 555 113 561 131
rect 579 113 585 131
rect 555 100 585 113
<< pdiffc >>
rect 121 869 139 887
rect 121 833 139 851
rect 121 797 139 815
rect 121 761 139 779
rect 121 725 139 743
rect 121 689 139 707
rect 121 653 139 671
rect 121 617 139 635
rect 121 581 139 599
rect 121 545 139 563
rect 121 509 139 527
rect 121 473 139 491
rect 121 437 139 455
rect 121 401 139 419
rect 121 365 139 383
rect 121 329 139 347
rect 121 293 139 311
rect 121 257 139 275
rect 121 221 139 239
rect 121 185 139 203
rect 121 149 139 167
rect 121 113 139 131
rect 341 869 359 887
rect 341 833 359 851
rect 341 797 359 815
rect 341 761 359 779
rect 341 725 359 743
rect 341 689 359 707
rect 341 653 359 671
rect 341 617 359 635
rect 341 581 359 599
rect 341 545 359 563
rect 341 509 359 527
rect 341 473 359 491
rect 341 437 359 455
rect 341 401 359 419
rect 341 365 359 383
rect 341 329 359 347
rect 341 293 359 311
rect 341 257 359 275
rect 341 221 359 239
rect 341 185 359 203
rect 341 149 359 167
rect 341 113 359 131
rect 561 869 579 887
rect 561 833 579 851
rect 561 797 579 815
rect 561 761 579 779
rect 561 725 579 743
rect 561 689 579 707
rect 561 653 579 671
rect 561 617 579 635
rect 561 581 579 599
rect 561 545 579 563
rect 561 509 579 527
rect 561 473 579 491
rect 561 437 579 455
rect 561 401 579 419
rect 561 365 579 383
rect 561 329 579 347
rect 561 293 579 311
rect 561 257 579 275
rect 561 221 579 239
rect 561 185 579 203
rect 561 149 579 167
rect 561 113 579 131
<< nsubdiff >>
rect 67 934 89 952
rect 107 934 125 952
rect 143 934 161 952
rect 179 934 197 952
rect 215 934 233 952
rect 251 934 269 952
rect 287 934 305 952
rect 323 934 341 952
rect 359 934 377 952
rect 395 934 413 952
rect 431 934 449 952
rect 467 934 485 952
rect 503 934 521 952
rect 539 934 557 952
rect 575 934 593 952
rect 611 934 633 952
rect 67 917 85 934
rect 615 917 633 934
rect 67 881 85 899
rect 67 845 85 863
rect 67 809 85 827
rect 67 773 85 791
rect 67 737 85 755
rect 67 701 85 719
rect 67 665 85 683
rect 67 629 85 647
rect 67 593 85 611
rect 67 557 85 575
rect 67 521 85 539
rect 67 485 85 503
rect 67 449 85 467
rect 67 413 85 431
rect 67 377 85 395
rect 67 341 85 359
rect 67 305 85 323
rect 67 269 85 287
rect 67 239 85 251
rect 615 881 633 899
rect 615 845 633 863
rect 615 809 633 827
rect 615 773 633 791
rect 615 737 633 755
rect 615 701 633 719
rect 615 665 633 683
rect 615 629 633 647
rect 615 593 633 611
rect 615 557 633 575
rect 615 521 633 539
rect 615 485 633 503
rect 615 449 633 467
rect 615 413 633 431
rect 615 377 633 395
rect 615 341 633 359
rect 615 305 633 323
rect 615 269 633 287
rect 615 239 633 251
<< nsubdiffcont >>
rect 89 934 107 952
rect 125 934 143 952
rect 161 934 179 952
rect 197 934 215 952
rect 233 934 251 952
rect 269 934 287 952
rect 305 934 323 952
rect 341 934 359 952
rect 377 934 395 952
rect 413 934 431 952
rect 449 934 467 952
rect 485 934 503 952
rect 521 934 539 952
rect 557 934 575 952
rect 593 934 611 952
rect 67 899 85 917
rect 67 863 85 881
rect 67 827 85 845
rect 67 791 85 809
rect 67 755 85 773
rect 67 719 85 737
rect 67 683 85 701
rect 67 647 85 665
rect 67 611 85 629
rect 67 575 85 593
rect 67 539 85 557
rect 67 503 85 521
rect 67 467 85 485
rect 67 431 85 449
rect 67 395 85 413
rect 67 359 85 377
rect 67 323 85 341
rect 67 287 85 305
rect 67 251 85 269
rect 615 899 633 917
rect 615 863 633 881
rect 615 827 633 845
rect 615 791 633 809
rect 615 755 633 773
rect 615 719 633 737
rect 615 683 633 701
rect 615 647 633 665
rect 615 611 633 629
rect 615 575 633 593
rect 615 539 633 557
rect 615 503 633 521
rect 615 467 633 485
rect 615 431 633 449
rect 615 395 633 413
rect 615 359 633 377
rect 615 323 633 341
rect 615 287 633 305
rect 615 251 633 269
<< poly >>
rect 145 900 335 913
rect 365 900 555 913
rect 145 50 335 100
rect 365 50 555 100
<< locali >>
rect 67 934 89 952
rect 107 934 125 952
rect 143 934 161 952
rect 179 934 197 952
rect 215 934 233 952
rect 251 934 269 952
rect 287 934 305 952
rect 323 934 341 952
rect 359 934 377 952
rect 395 934 413 952
rect 431 934 449 952
rect 467 934 485 952
rect 503 934 521 952
rect 539 934 557 952
rect 575 934 593 952
rect 611 934 633 952
rect 67 917 85 934
rect 67 881 85 899
rect 67 845 85 863
rect 67 809 85 827
rect 67 773 85 791
rect 67 737 85 755
rect 67 701 85 719
rect 67 665 85 683
rect 67 629 85 647
rect 67 593 85 611
rect 67 557 85 575
rect 67 521 85 539
rect 67 485 85 503
rect 67 449 85 467
rect 67 413 85 431
rect 67 377 85 395
rect 67 341 85 359
rect 67 305 85 323
rect 67 269 85 287
rect 67 239 85 251
rect 115 887 145 934
rect 115 869 121 887
rect 139 869 145 887
rect 115 851 145 869
rect 115 833 121 851
rect 139 833 145 851
rect 115 815 145 833
rect 115 797 121 815
rect 139 797 145 815
rect 115 779 145 797
rect 115 761 121 779
rect 139 761 145 779
rect 115 743 145 761
rect 115 725 121 743
rect 139 725 145 743
rect 115 707 145 725
rect 115 689 121 707
rect 139 689 145 707
rect 115 671 145 689
rect 115 653 121 671
rect 139 653 145 671
rect 115 635 145 653
rect 115 617 121 635
rect 139 617 145 635
rect 115 599 145 617
rect 115 581 121 599
rect 139 581 145 599
rect 115 563 145 581
rect 115 545 121 563
rect 139 545 145 563
rect 115 527 145 545
rect 115 509 121 527
rect 139 509 145 527
rect 115 491 145 509
rect 115 473 121 491
rect 139 473 145 491
rect 115 455 145 473
rect 115 437 121 455
rect 139 437 145 455
rect 115 419 145 437
rect 115 401 121 419
rect 139 401 145 419
rect 115 383 145 401
rect 115 365 121 383
rect 139 365 145 383
rect 115 347 145 365
rect 115 329 121 347
rect 139 329 145 347
rect 115 311 145 329
rect 115 293 121 311
rect 139 293 145 311
rect 115 275 145 293
rect 115 257 121 275
rect 139 257 145 275
rect 115 239 145 257
rect 115 221 121 239
rect 139 221 145 239
rect 115 203 145 221
rect 115 185 121 203
rect 139 185 145 203
rect 115 167 145 185
rect 115 149 121 167
rect 139 149 145 167
rect 115 131 145 149
rect 115 113 121 131
rect 139 113 145 131
rect 115 98 145 113
rect 335 887 365 902
rect 335 869 341 887
rect 359 869 365 887
rect 335 851 365 869
rect 335 833 341 851
rect 359 833 365 851
rect 335 815 365 833
rect 335 797 341 815
rect 359 797 365 815
rect 335 779 365 797
rect 335 761 341 779
rect 359 761 365 779
rect 335 743 365 761
rect 335 725 341 743
rect 359 725 365 743
rect 335 707 365 725
rect 335 689 341 707
rect 359 689 365 707
rect 335 671 365 689
rect 335 653 341 671
rect 359 653 365 671
rect 335 635 365 653
rect 335 617 341 635
rect 359 617 365 635
rect 335 599 365 617
rect 335 581 341 599
rect 359 581 365 599
rect 335 563 365 581
rect 335 545 341 563
rect 359 545 365 563
rect 335 527 365 545
rect 335 509 341 527
rect 359 509 365 527
rect 335 491 365 509
rect 335 473 341 491
rect 359 473 365 491
rect 335 455 365 473
rect 335 437 341 455
rect 359 437 365 455
rect 335 419 365 437
rect 335 401 341 419
rect 359 401 365 419
rect 335 383 365 401
rect 335 365 341 383
rect 359 365 365 383
rect 335 347 365 365
rect 335 329 341 347
rect 359 329 365 347
rect 335 311 365 329
rect 335 293 341 311
rect 359 293 365 311
rect 335 275 365 293
rect 335 257 341 275
rect 359 257 365 275
rect 335 239 365 257
rect 335 221 341 239
rect 359 221 365 239
rect 335 203 365 221
rect 335 185 341 203
rect 359 185 365 203
rect 335 167 365 185
rect 335 149 341 167
rect 359 149 365 167
rect 335 131 365 149
rect 335 113 341 131
rect 359 113 365 131
rect 335 98 365 113
rect 555 887 585 934
rect 555 869 561 887
rect 579 869 585 887
rect 555 851 585 869
rect 555 833 561 851
rect 579 833 585 851
rect 555 815 585 833
rect 555 797 561 815
rect 579 797 585 815
rect 555 779 585 797
rect 555 761 561 779
rect 579 761 585 779
rect 555 743 585 761
rect 555 725 561 743
rect 579 725 585 743
rect 555 707 585 725
rect 555 689 561 707
rect 579 689 585 707
rect 555 671 585 689
rect 555 653 561 671
rect 579 653 585 671
rect 555 635 585 653
rect 555 617 561 635
rect 579 617 585 635
rect 555 599 585 617
rect 555 581 561 599
rect 579 581 585 599
rect 555 563 585 581
rect 555 545 561 563
rect 579 545 585 563
rect 555 527 585 545
rect 555 509 561 527
rect 579 509 585 527
rect 555 491 585 509
rect 555 473 561 491
rect 579 473 585 491
rect 555 455 585 473
rect 555 437 561 455
rect 579 437 585 455
rect 555 419 585 437
rect 555 401 561 419
rect 579 401 585 419
rect 555 383 585 401
rect 555 365 561 383
rect 579 365 585 383
rect 555 347 585 365
rect 555 329 561 347
rect 579 329 585 347
rect 555 311 585 329
rect 555 293 561 311
rect 579 293 585 311
rect 555 275 585 293
rect 555 257 561 275
rect 579 257 585 275
rect 555 239 585 257
rect 615 917 633 934
rect 615 881 633 899
rect 615 845 633 863
rect 615 809 633 827
rect 615 773 633 791
rect 615 737 633 755
rect 615 701 633 719
rect 615 665 633 683
rect 615 629 633 647
rect 615 593 633 611
rect 615 557 633 575
rect 615 521 633 539
rect 615 485 633 503
rect 615 449 633 467
rect 615 413 633 431
rect 615 377 633 395
rect 615 341 633 359
rect 615 305 633 323
rect 615 269 633 287
rect 615 239 633 251
rect 555 221 561 239
rect 579 221 585 239
rect 555 203 585 221
rect 555 185 561 203
rect 579 185 585 203
rect 555 167 585 185
rect 555 149 561 167
rect 579 149 585 167
rect 555 131 585 149
rect 555 113 561 131
rect 579 113 585 131
rect 555 98 585 113
<< end >>
