magic
tech sky130A
magscale 1 2
timestamp 1622803027
<< nwell >>
rect 100 1640 1270 2815
rect 3695 1752 4447 2814
rect 2266 537 3436 1708
rect 4990 547 5742 1602
<< pwell >>
rect 1430 2092 3436 3372
rect 4572 2349 5742 3371
rect 4571 2339 5742 2349
rect 4571 2151 5741 2339
rect 100 -10 2106 1202
rect 3695 -10 4865 1210
<< nmos >>
rect 1626 2302 1986 3202
rect 2044 2302 2404 3202
rect 2462 2302 2822 3202
rect 2880 2302 3240 3202
rect 4768 2399 5128 3199
rect 5186 2399 5546 3199
rect 296 160 656 1060
rect 714 160 1074 1060
rect 1132 160 1492 1060
rect 1550 160 1910 1060
rect 3891 162 4251 962
rect 4309 162 4669 962
<< pmos >>
rect 296 1754 656 2654
rect 714 1754 1074 2654
rect 3891 1843 4251 2643
rect 2462 698 2822 1598
rect 2880 698 3240 1598
rect 5186 718 5546 1518
<< ndiff >>
rect 1568 3190 1626 3202
rect 1568 3140 1580 3190
rect 1614 3140 1626 3190
rect 1568 3100 1626 3140
rect 1568 3060 1580 3100
rect 1614 3060 1626 3100
rect 1568 3020 1626 3060
rect 1568 2980 1580 3020
rect 1614 2980 1626 3020
rect 1568 2940 1626 2980
rect 1568 2900 1580 2940
rect 1614 2900 1626 2940
rect 1568 2860 1626 2900
rect 1568 2820 1580 2860
rect 1614 2820 1626 2860
rect 1568 2780 1626 2820
rect 1568 2740 1580 2780
rect 1614 2740 1626 2780
rect 1568 2700 1626 2740
rect 1568 2660 1580 2700
rect 1614 2660 1626 2700
rect 1568 2620 1626 2660
rect 1568 2580 1580 2620
rect 1614 2580 1626 2620
rect 1568 2540 1626 2580
rect 1568 2500 1580 2540
rect 1614 2500 1626 2540
rect 1568 2460 1626 2500
rect 1568 2420 1580 2460
rect 1614 2420 1626 2460
rect 1568 2380 1626 2420
rect 1568 2314 1580 2380
rect 1614 2314 1626 2380
rect 1568 2302 1626 2314
rect 1986 3190 2044 3202
rect 1986 3140 1998 3190
rect 2032 3140 2044 3190
rect 1986 3100 2044 3140
rect 1986 3060 1998 3100
rect 2032 3060 2044 3100
rect 1986 3020 2044 3060
rect 1986 2980 1998 3020
rect 2032 2980 2044 3020
rect 1986 2940 2044 2980
rect 1986 2900 1998 2940
rect 2032 2900 2044 2940
rect 1986 2860 2044 2900
rect 1986 2820 1998 2860
rect 2032 2820 2044 2860
rect 1986 2780 2044 2820
rect 1986 2740 1998 2780
rect 2032 2740 2044 2780
rect 1986 2700 2044 2740
rect 1986 2660 1998 2700
rect 2032 2660 2044 2700
rect 1986 2620 2044 2660
rect 1986 2580 1998 2620
rect 2032 2580 2044 2620
rect 1986 2540 2044 2580
rect 1986 2500 1998 2540
rect 2032 2500 2044 2540
rect 1986 2460 2044 2500
rect 1986 2420 1998 2460
rect 2032 2420 2044 2460
rect 1986 2380 2044 2420
rect 1986 2314 1998 2380
rect 2032 2314 2044 2380
rect 1986 2302 2044 2314
rect 2404 3190 2462 3202
rect 2404 3140 2416 3190
rect 2450 3140 2462 3190
rect 2404 3100 2462 3140
rect 2404 3060 2416 3100
rect 2450 3060 2462 3100
rect 2404 3020 2462 3060
rect 2404 2980 2416 3020
rect 2450 2980 2462 3020
rect 2404 2940 2462 2980
rect 2404 2900 2416 2940
rect 2450 2900 2462 2940
rect 2404 2860 2462 2900
rect 2404 2820 2416 2860
rect 2450 2820 2462 2860
rect 2404 2780 2462 2820
rect 2404 2740 2416 2780
rect 2450 2740 2462 2780
rect 2404 2700 2462 2740
rect 2404 2660 2416 2700
rect 2450 2660 2462 2700
rect 2404 2620 2462 2660
rect 2404 2580 2416 2620
rect 2450 2580 2462 2620
rect 2404 2540 2462 2580
rect 2404 2500 2416 2540
rect 2450 2500 2462 2540
rect 2404 2460 2462 2500
rect 2404 2420 2416 2460
rect 2450 2420 2462 2460
rect 2404 2380 2462 2420
rect 2404 2340 2416 2380
rect 2450 2340 2462 2380
rect 2404 2302 2462 2340
rect 2822 3190 2880 3202
rect 2822 3152 2834 3190
rect 2868 3152 2880 3190
rect 2822 3112 2880 3152
rect 2822 3072 2834 3112
rect 2868 3072 2880 3112
rect 2822 3032 2880 3072
rect 2822 2992 2834 3032
rect 2868 2992 2880 3032
rect 2822 2952 2880 2992
rect 2822 2912 2834 2952
rect 2868 2912 2880 2952
rect 2822 2872 2880 2912
rect 2822 2832 2834 2872
rect 2868 2832 2880 2872
rect 2822 2792 2880 2832
rect 2822 2752 2834 2792
rect 2868 2752 2880 2792
rect 2822 2712 2880 2752
rect 2822 2672 2834 2712
rect 2868 2672 2880 2712
rect 2822 2632 2880 2672
rect 2822 2592 2834 2632
rect 2868 2592 2880 2632
rect 2822 2552 2880 2592
rect 2822 2512 2834 2552
rect 2868 2512 2880 2552
rect 2822 2472 2880 2512
rect 2822 2432 2834 2472
rect 2868 2432 2880 2472
rect 2822 2392 2880 2432
rect 2822 2352 2834 2392
rect 2868 2352 2880 2392
rect 2822 2302 2880 2352
rect 3240 3190 3298 3202
rect 3240 3140 3252 3190
rect 3286 3140 3298 3190
rect 3240 3100 3298 3140
rect 3240 3060 3252 3100
rect 3286 3060 3298 3100
rect 3240 3020 3298 3060
rect 3240 2980 3252 3020
rect 3286 2980 3298 3020
rect 3240 2940 3298 2980
rect 3240 2900 3252 2940
rect 3286 2900 3298 2940
rect 3240 2860 3298 2900
rect 3240 2820 3252 2860
rect 3286 2820 3298 2860
rect 3240 2780 3298 2820
rect 3240 2740 3252 2780
rect 3286 2740 3298 2780
rect 4710 3187 4768 3199
rect 4710 3139 4722 3187
rect 4756 3139 4768 3187
rect 4710 3099 4768 3139
rect 4710 3059 4722 3099
rect 4756 3059 4768 3099
rect 4710 3019 4768 3059
rect 4710 2979 4722 3019
rect 4756 2979 4768 3019
rect 4710 2939 4768 2979
rect 4710 2899 4722 2939
rect 4756 2899 4768 2939
rect 4710 2859 4768 2899
rect 4710 2819 4722 2859
rect 4756 2819 4768 2859
rect 4710 2779 4768 2819
rect 3240 2700 3298 2740
rect 3240 2660 3252 2700
rect 3286 2660 3298 2700
rect 3240 2620 3298 2660
rect 3240 2580 3252 2620
rect 3286 2580 3298 2620
rect 3240 2540 3298 2580
rect 3240 2500 3252 2540
rect 3286 2500 3298 2540
rect 3240 2460 3298 2500
rect 3240 2420 3252 2460
rect 3286 2420 3298 2460
rect 3240 2380 3298 2420
rect 3240 2340 3252 2380
rect 3286 2340 3298 2380
rect 3240 2302 3298 2340
rect 4710 2739 4722 2779
rect 4756 2739 4768 2779
rect 4710 2699 4768 2739
rect 4710 2659 4722 2699
rect 4756 2659 4768 2699
rect 4710 2619 4768 2659
rect 4710 2579 4722 2619
rect 4756 2579 4768 2619
rect 4710 2539 4768 2579
rect 4710 2499 4722 2539
rect 4756 2499 4768 2539
rect 4710 2459 4768 2499
rect 4710 2411 4722 2459
rect 4756 2411 4768 2459
rect 4710 2399 4768 2411
rect 5128 3187 5186 3199
rect 5128 3139 5140 3187
rect 5174 3139 5186 3187
rect 5128 3099 5186 3139
rect 5128 3059 5140 3099
rect 5174 3059 5186 3099
rect 5128 3019 5186 3059
rect 5128 2979 5140 3019
rect 5174 2979 5186 3019
rect 5128 2939 5186 2979
rect 5128 2899 5140 2939
rect 5174 2899 5186 2939
rect 5128 2859 5186 2899
rect 5128 2819 5140 2859
rect 5174 2819 5186 2859
rect 5128 2779 5186 2819
rect 5128 2739 5140 2779
rect 5174 2739 5186 2779
rect 5128 2699 5186 2739
rect 5128 2659 5140 2699
rect 5174 2659 5186 2699
rect 5128 2619 5186 2659
rect 5128 2579 5140 2619
rect 5174 2579 5186 2619
rect 5128 2539 5186 2579
rect 5128 2499 5140 2539
rect 5174 2499 5186 2539
rect 5128 2459 5186 2499
rect 5128 2411 5140 2459
rect 5174 2411 5186 2459
rect 5128 2399 5186 2411
rect 5546 3187 5604 3199
rect 5546 3139 5558 3187
rect 5592 3139 5604 3187
rect 5546 3099 5604 3139
rect 5546 3059 5558 3099
rect 5592 3059 5604 3099
rect 5546 3019 5604 3059
rect 5546 2979 5558 3019
rect 5592 2979 5604 3019
rect 5546 2939 5604 2979
rect 5546 2899 5558 2939
rect 5592 2899 5604 2939
rect 5546 2859 5604 2899
rect 5546 2819 5558 2859
rect 5592 2819 5604 2859
rect 5546 2779 5604 2819
rect 5546 2739 5558 2779
rect 5592 2739 5604 2779
rect 5546 2699 5604 2739
rect 5546 2659 5558 2699
rect 5592 2659 5604 2699
rect 5546 2619 5604 2659
rect 5546 2579 5558 2619
rect 5592 2579 5604 2619
rect 5546 2539 5604 2579
rect 5546 2499 5558 2539
rect 5592 2499 5604 2539
rect 5546 2459 5604 2499
rect 5546 2411 5558 2459
rect 5592 2411 5604 2459
rect 5546 2399 5604 2411
rect 238 1022 296 1060
rect 238 982 250 1022
rect 284 982 296 1022
rect 238 942 296 982
rect 238 902 250 942
rect 284 902 296 942
rect 238 862 296 902
rect 238 822 250 862
rect 284 822 296 862
rect 238 782 296 822
rect 238 742 250 782
rect 284 742 296 782
rect 238 702 296 742
rect 238 662 250 702
rect 284 662 296 702
rect 238 622 296 662
rect 238 582 250 622
rect 284 582 296 622
rect 238 542 296 582
rect 238 502 250 542
rect 284 502 296 542
rect 238 462 296 502
rect 238 422 250 462
rect 284 422 296 462
rect 238 382 296 422
rect 238 342 250 382
rect 284 342 296 382
rect 238 302 296 342
rect 238 262 250 302
rect 284 262 296 302
rect 238 222 296 262
rect 238 172 250 222
rect 284 172 296 222
rect 238 160 296 172
rect 656 1010 714 1060
rect 656 970 668 1010
rect 702 970 714 1010
rect 656 930 714 970
rect 656 890 668 930
rect 702 890 714 930
rect 656 850 714 890
rect 656 810 668 850
rect 702 810 714 850
rect 656 770 714 810
rect 656 730 668 770
rect 702 730 714 770
rect 656 690 714 730
rect 656 650 668 690
rect 702 650 714 690
rect 656 610 714 650
rect 656 570 668 610
rect 702 570 714 610
rect 656 530 714 570
rect 656 490 668 530
rect 702 490 714 530
rect 656 450 714 490
rect 656 410 668 450
rect 702 410 714 450
rect 656 370 714 410
rect 656 330 668 370
rect 702 330 714 370
rect 656 290 714 330
rect 656 250 668 290
rect 702 250 714 290
rect 656 210 714 250
rect 656 172 668 210
rect 702 172 714 210
rect 656 160 714 172
rect 1074 1022 1132 1060
rect 1074 982 1086 1022
rect 1120 982 1132 1022
rect 1074 942 1132 982
rect 1074 902 1086 942
rect 1120 902 1132 942
rect 1074 862 1132 902
rect 1074 822 1086 862
rect 1120 822 1132 862
rect 1074 782 1132 822
rect 1074 742 1086 782
rect 1120 742 1132 782
rect 1074 702 1132 742
rect 1074 662 1086 702
rect 1120 662 1132 702
rect 1074 622 1132 662
rect 1074 582 1086 622
rect 1120 582 1132 622
rect 1074 542 1132 582
rect 1074 502 1086 542
rect 1120 502 1132 542
rect 1074 462 1132 502
rect 1074 422 1086 462
rect 1120 422 1132 462
rect 1074 382 1132 422
rect 1074 342 1086 382
rect 1120 342 1132 382
rect 1074 302 1132 342
rect 1074 262 1086 302
rect 1120 262 1132 302
rect 1074 222 1132 262
rect 1074 172 1086 222
rect 1120 172 1132 222
rect 1074 160 1132 172
rect 1492 1048 1550 1060
rect 1492 982 1504 1048
rect 1538 982 1550 1048
rect 1492 942 1550 982
rect 1492 902 1504 942
rect 1538 902 1550 942
rect 1492 862 1550 902
rect 1492 822 1504 862
rect 1538 822 1550 862
rect 1492 782 1550 822
rect 1492 742 1504 782
rect 1538 742 1550 782
rect 1492 702 1550 742
rect 1492 662 1504 702
rect 1538 662 1550 702
rect 1492 622 1550 662
rect 1492 582 1504 622
rect 1538 582 1550 622
rect 1492 542 1550 582
rect 1492 502 1504 542
rect 1538 502 1550 542
rect 1492 462 1550 502
rect 1492 422 1504 462
rect 1538 422 1550 462
rect 1492 382 1550 422
rect 1492 342 1504 382
rect 1538 342 1550 382
rect 1492 302 1550 342
rect 1492 262 1504 302
rect 1538 262 1550 302
rect 1492 222 1550 262
rect 1492 172 1504 222
rect 1538 172 1550 222
rect 1492 160 1550 172
rect 1910 1048 1968 1060
rect 1910 982 1922 1048
rect 1956 982 1968 1048
rect 1910 942 1968 982
rect 1910 902 1922 942
rect 1956 902 1968 942
rect 1910 862 1968 902
rect 1910 822 1922 862
rect 1956 822 1968 862
rect 1910 782 1968 822
rect 1910 742 1922 782
rect 1956 742 1968 782
rect 1910 702 1968 742
rect 1910 662 1922 702
rect 1956 662 1968 702
rect 1910 622 1968 662
rect 1910 582 1922 622
rect 1956 582 1968 622
rect 1910 542 1968 582
rect 3833 950 3891 962
rect 3833 902 3845 950
rect 3879 902 3891 950
rect 3833 862 3891 902
rect 3833 822 3845 862
rect 3879 822 3891 862
rect 3833 782 3891 822
rect 3833 742 3845 782
rect 3879 742 3891 782
rect 3833 702 3891 742
rect 3833 662 3845 702
rect 3879 662 3891 702
rect 3833 622 3891 662
rect 3833 582 3845 622
rect 3879 582 3891 622
rect 1910 502 1922 542
rect 1956 502 1968 542
rect 1910 462 1968 502
rect 1910 422 1922 462
rect 1956 422 1968 462
rect 1910 382 1968 422
rect 1910 342 1922 382
rect 1956 342 1968 382
rect 1910 302 1968 342
rect 1910 262 1922 302
rect 1956 262 1968 302
rect 1910 222 1968 262
rect 1910 172 1922 222
rect 1956 172 1968 222
rect 1910 160 1968 172
rect 3833 542 3891 582
rect 3833 502 3845 542
rect 3879 502 3891 542
rect 3833 462 3891 502
rect 3833 422 3845 462
rect 3879 422 3891 462
rect 3833 382 3891 422
rect 3833 342 3845 382
rect 3879 342 3891 382
rect 3833 302 3891 342
rect 3833 262 3845 302
rect 3879 262 3891 302
rect 3833 222 3891 262
rect 3833 174 3845 222
rect 3879 174 3891 222
rect 3833 162 3891 174
rect 4251 950 4309 962
rect 4251 902 4263 950
rect 4297 902 4309 950
rect 4251 862 4309 902
rect 4251 822 4263 862
rect 4297 822 4309 862
rect 4251 782 4309 822
rect 4251 742 4263 782
rect 4297 742 4309 782
rect 4251 702 4309 742
rect 4251 662 4263 702
rect 4297 662 4309 702
rect 4251 622 4309 662
rect 4251 582 4263 622
rect 4297 582 4309 622
rect 4251 542 4309 582
rect 4251 502 4263 542
rect 4297 502 4309 542
rect 4251 462 4309 502
rect 4251 422 4263 462
rect 4297 422 4309 462
rect 4251 382 4309 422
rect 4251 342 4263 382
rect 4297 342 4309 382
rect 4251 302 4309 342
rect 4251 262 4263 302
rect 4297 262 4309 302
rect 4251 222 4309 262
rect 4251 174 4263 222
rect 4297 174 4309 222
rect 4251 162 4309 174
rect 4669 950 4727 962
rect 4669 902 4681 950
rect 4715 902 4727 950
rect 4669 862 4727 902
rect 4669 822 4681 862
rect 4715 822 4727 862
rect 4669 782 4727 822
rect 4669 742 4681 782
rect 4715 742 4727 782
rect 4669 702 4727 742
rect 4669 662 4681 702
rect 4715 662 4727 702
rect 4669 622 4727 662
rect 4669 582 4681 622
rect 4715 582 4727 622
rect 4669 542 4727 582
rect 4669 502 4681 542
rect 4715 502 4727 542
rect 4669 462 4727 502
rect 4669 422 4681 462
rect 4715 422 4727 462
rect 4669 382 4727 422
rect 4669 342 4681 382
rect 4715 342 4727 382
rect 4669 302 4727 342
rect 4669 262 4681 302
rect 4715 262 4727 302
rect 4669 222 4727 262
rect 4669 174 4681 222
rect 4715 174 4727 222
rect 4669 162 4727 174
<< pdiff >>
rect 238 2642 296 2654
rect 238 2600 250 2642
rect 284 2600 296 2642
rect 238 2560 296 2600
rect 238 2520 250 2560
rect 284 2520 296 2560
rect 238 2480 296 2520
rect 238 2440 250 2480
rect 284 2440 296 2480
rect 238 2400 296 2440
rect 238 2360 250 2400
rect 284 2360 296 2400
rect 238 2320 296 2360
rect 238 2280 250 2320
rect 284 2280 296 2320
rect 238 2240 296 2280
rect 238 2200 250 2240
rect 284 2200 296 2240
rect 238 2160 296 2200
rect 238 2120 250 2160
rect 284 2120 296 2160
rect 238 2080 296 2120
rect 238 2040 250 2080
rect 284 2040 296 2080
rect 238 2000 296 2040
rect 238 1960 250 2000
rect 284 1960 296 2000
rect 238 1920 296 1960
rect 238 1880 250 1920
rect 284 1880 296 1920
rect 238 1840 296 1880
rect 238 1800 250 1840
rect 284 1800 296 1840
rect 238 1754 296 1800
rect 656 2608 714 2654
rect 656 2568 668 2608
rect 702 2568 714 2608
rect 656 2528 714 2568
rect 656 2488 668 2528
rect 702 2488 714 2528
rect 656 2448 714 2488
rect 656 2408 668 2448
rect 702 2408 714 2448
rect 656 2368 714 2408
rect 656 2328 668 2368
rect 702 2328 714 2368
rect 656 2288 714 2328
rect 656 2248 668 2288
rect 702 2248 714 2288
rect 656 2208 714 2248
rect 656 2168 668 2208
rect 702 2168 714 2208
rect 656 2128 714 2168
rect 656 2088 668 2128
rect 702 2088 714 2128
rect 656 2048 714 2088
rect 656 2008 668 2048
rect 702 2008 714 2048
rect 656 1968 714 2008
rect 656 1928 668 1968
rect 702 1928 714 1968
rect 656 1888 714 1928
rect 656 1848 668 1888
rect 702 1848 714 1888
rect 656 1808 714 1848
rect 656 1766 668 1808
rect 702 1766 714 1808
rect 656 1754 714 1766
rect 1074 2642 1132 2654
rect 1074 2600 1086 2642
rect 1120 2600 1132 2642
rect 1074 2560 1132 2600
rect 1074 2520 1086 2560
rect 1120 2520 1132 2560
rect 1074 2480 1132 2520
rect 1074 2440 1086 2480
rect 1120 2440 1132 2480
rect 1074 2400 1132 2440
rect 1074 2360 1086 2400
rect 1120 2360 1132 2400
rect 1074 2320 1132 2360
rect 1074 2280 1086 2320
rect 1120 2280 1132 2320
rect 1074 2240 1132 2280
rect 1074 2200 1086 2240
rect 1120 2200 1132 2240
rect 1074 2160 1132 2200
rect 1074 2120 1086 2160
rect 1120 2120 1132 2160
rect 1074 2080 1132 2120
rect 1074 2040 1086 2080
rect 1120 2040 1132 2080
rect 1074 2000 1132 2040
rect 1074 1960 1086 2000
rect 1120 1960 1132 2000
rect 1074 1920 1132 1960
rect 1074 1880 1086 1920
rect 1120 1880 1132 1920
rect 1074 1840 1132 1880
rect 1074 1800 1086 1840
rect 1120 1800 1132 1840
rect 1074 1754 1132 1800
rect 3833 2631 3891 2643
rect 3833 2580 3845 2631
rect 3879 2580 3891 2631
rect 3833 2540 3891 2580
rect 3833 2500 3845 2540
rect 3879 2500 3891 2540
rect 3833 2460 3891 2500
rect 3833 2420 3845 2460
rect 3879 2420 3891 2460
rect 3833 2380 3891 2420
rect 3833 2340 3845 2380
rect 3879 2340 3891 2380
rect 3833 2300 3891 2340
rect 3833 2260 3845 2300
rect 3879 2260 3891 2300
rect 3833 2220 3891 2260
rect 3833 2180 3845 2220
rect 3879 2180 3891 2220
rect 3833 2140 3891 2180
rect 3833 2100 3845 2140
rect 3879 2100 3891 2140
rect 3833 2060 3891 2100
rect 3833 2020 3845 2060
rect 3879 2020 3891 2060
rect 3833 1980 3891 2020
rect 3833 1922 3845 1980
rect 3879 1922 3891 1980
rect 3833 1843 3891 1922
rect 4251 2631 4309 2643
rect 4251 2580 4263 2631
rect 4297 2580 4309 2631
rect 4251 2540 4309 2580
rect 4251 2500 4263 2540
rect 4297 2500 4309 2540
rect 4251 2460 4309 2500
rect 4251 2420 4263 2460
rect 4297 2420 4309 2460
rect 4251 2380 4309 2420
rect 4251 2340 4263 2380
rect 4297 2340 4309 2380
rect 4251 2300 4309 2340
rect 4251 2260 4263 2300
rect 4297 2260 4309 2300
rect 4251 2220 4309 2260
rect 4251 2180 4263 2220
rect 4297 2180 4309 2220
rect 4251 2140 4309 2180
rect 4251 2100 4263 2140
rect 4297 2100 4309 2140
rect 4251 2060 4309 2100
rect 4251 2020 4263 2060
rect 4297 2020 4309 2060
rect 4251 1980 4309 2020
rect 4251 1940 4263 1980
rect 4297 1940 4309 1980
rect 4251 1900 4309 1940
rect 4251 1855 4263 1900
rect 4297 1855 4309 1900
rect 4251 1843 4309 1855
rect 2404 1552 2462 1598
rect 2404 1512 2416 1552
rect 2450 1512 2462 1552
rect 2404 1472 2462 1512
rect 2404 1432 2416 1472
rect 2450 1432 2462 1472
rect 2404 1392 2462 1432
rect 2404 1352 2416 1392
rect 2450 1352 2462 1392
rect 2404 1312 2462 1352
rect 2404 1272 2416 1312
rect 2450 1272 2462 1312
rect 2404 1232 2462 1272
rect 2404 1192 2416 1232
rect 2450 1192 2462 1232
rect 2404 1152 2462 1192
rect 2404 1112 2416 1152
rect 2450 1112 2462 1152
rect 2404 1072 2462 1112
rect 2404 1032 2416 1072
rect 2450 1032 2462 1072
rect 2404 992 2462 1032
rect 2404 952 2416 992
rect 2450 952 2462 992
rect 2404 912 2462 952
rect 2404 872 2416 912
rect 2450 872 2462 912
rect 2404 832 2462 872
rect 2404 792 2416 832
rect 2450 792 2462 832
rect 2404 752 2462 792
rect 2404 710 2416 752
rect 2450 710 2462 752
rect 2404 698 2462 710
rect 2822 1586 2880 1598
rect 2822 1544 2834 1586
rect 2868 1544 2880 1586
rect 2822 1504 2880 1544
rect 2822 1464 2834 1504
rect 2868 1464 2880 1504
rect 2822 1424 2880 1464
rect 2822 1384 2834 1424
rect 2868 1384 2880 1424
rect 2822 1344 2880 1384
rect 2822 1304 2834 1344
rect 2868 1304 2880 1344
rect 2822 1264 2880 1304
rect 2822 1224 2834 1264
rect 2868 1224 2880 1264
rect 2822 1184 2880 1224
rect 2822 1144 2834 1184
rect 2868 1144 2880 1184
rect 2822 1104 2880 1144
rect 2822 1064 2834 1104
rect 2868 1064 2880 1104
rect 2822 1024 2880 1064
rect 2822 984 2834 1024
rect 2868 984 2880 1024
rect 2822 944 2880 984
rect 2822 904 2834 944
rect 2868 904 2880 944
rect 2822 864 2880 904
rect 2822 824 2834 864
rect 2868 824 2880 864
rect 2822 784 2880 824
rect 2822 744 2834 784
rect 2868 744 2880 784
rect 2822 698 2880 744
rect 3240 1552 3298 1598
rect 3240 1512 3252 1552
rect 3286 1512 3298 1552
rect 3240 1472 3298 1512
rect 3240 1432 3252 1472
rect 3286 1432 3298 1472
rect 3240 1392 3298 1432
rect 3240 1352 3252 1392
rect 3286 1352 3298 1392
rect 3240 1312 3298 1352
rect 3240 1272 3252 1312
rect 3286 1272 3298 1312
rect 3240 1232 3298 1272
rect 3240 1192 3252 1232
rect 3286 1192 3298 1232
rect 3240 1152 3298 1192
rect 3240 1112 3252 1152
rect 3286 1112 3298 1152
rect 3240 1072 3298 1112
rect 3240 1032 3252 1072
rect 3286 1032 3298 1072
rect 3240 992 3298 1032
rect 3240 952 3252 992
rect 3286 952 3298 992
rect 3240 912 3298 952
rect 3240 872 3252 912
rect 3286 872 3298 912
rect 3240 832 3298 872
rect 3240 792 3252 832
rect 3286 792 3298 832
rect 3240 752 3298 792
rect 3240 710 3252 752
rect 3286 710 3298 752
rect 3240 698 3298 710
rect 5128 1506 5186 1518
rect 5128 1462 5140 1506
rect 5174 1462 5186 1506
rect 5128 1422 5186 1462
rect 5128 1382 5140 1422
rect 5174 1382 5186 1422
rect 5128 1342 5186 1382
rect 5128 1302 5140 1342
rect 5174 1302 5186 1342
rect 5128 1262 5186 1302
rect 5128 1222 5140 1262
rect 5174 1222 5186 1262
rect 5128 1182 5186 1222
rect 5128 1142 5140 1182
rect 5174 1142 5186 1182
rect 5128 1102 5186 1142
rect 5128 1062 5140 1102
rect 5174 1062 5186 1102
rect 5128 1022 5186 1062
rect 5128 982 5140 1022
rect 5174 982 5186 1022
rect 5128 942 5186 982
rect 5128 902 5140 942
rect 5174 902 5186 942
rect 5128 862 5186 902
rect 5128 822 5140 862
rect 5174 822 5186 862
rect 5128 782 5186 822
rect 5128 730 5140 782
rect 5174 730 5186 782
rect 5128 718 5186 730
rect 5546 1506 5604 1518
rect 5546 1462 5558 1506
rect 5592 1462 5604 1506
rect 5546 1422 5604 1462
rect 5546 1382 5558 1422
rect 5592 1382 5604 1422
rect 5546 1342 5604 1382
rect 5546 1302 5558 1342
rect 5592 1302 5604 1342
rect 5546 1262 5604 1302
rect 5546 1222 5558 1262
rect 5592 1222 5604 1262
rect 5546 1182 5604 1222
rect 5546 1142 5558 1182
rect 5592 1142 5604 1182
rect 5546 1102 5604 1142
rect 5546 1062 5558 1102
rect 5592 1062 5604 1102
rect 5546 1022 5604 1062
rect 5546 982 5558 1022
rect 5592 982 5604 1022
rect 5546 942 5604 982
rect 5546 902 5558 942
rect 5592 902 5604 942
rect 5546 862 5604 902
rect 5546 822 5558 862
rect 5592 822 5604 862
rect 5546 782 5604 822
rect 5546 730 5558 782
rect 5592 730 5604 782
rect 5546 718 5604 730
<< ndiffc >>
rect 1580 3140 1614 3190
rect 1580 3060 1614 3100
rect 1580 2980 1614 3020
rect 1580 2900 1614 2940
rect 1580 2820 1614 2860
rect 1580 2740 1614 2780
rect 1580 2660 1614 2700
rect 1580 2580 1614 2620
rect 1580 2500 1614 2540
rect 1580 2420 1614 2460
rect 1580 2314 1614 2380
rect 1998 3140 2032 3190
rect 1998 3060 2032 3100
rect 1998 2980 2032 3020
rect 1998 2900 2032 2940
rect 1998 2820 2032 2860
rect 1998 2740 2032 2780
rect 1998 2660 2032 2700
rect 1998 2580 2032 2620
rect 1998 2500 2032 2540
rect 1998 2420 2032 2460
rect 1998 2314 2032 2380
rect 2416 3140 2450 3190
rect 2416 3060 2450 3100
rect 2416 2980 2450 3020
rect 2416 2900 2450 2940
rect 2416 2820 2450 2860
rect 2416 2740 2450 2780
rect 2416 2660 2450 2700
rect 2416 2580 2450 2620
rect 2416 2500 2450 2540
rect 2416 2420 2450 2460
rect 2416 2340 2450 2380
rect 2834 3152 2868 3190
rect 2834 3072 2868 3112
rect 2834 2992 2868 3032
rect 2834 2912 2868 2952
rect 2834 2832 2868 2872
rect 2834 2752 2868 2792
rect 2834 2672 2868 2712
rect 2834 2592 2868 2632
rect 2834 2512 2868 2552
rect 2834 2432 2868 2472
rect 2834 2352 2868 2392
rect 3252 3140 3286 3190
rect 3252 3060 3286 3100
rect 3252 2980 3286 3020
rect 3252 2900 3286 2940
rect 3252 2820 3286 2860
rect 3252 2740 3286 2780
rect 4722 3139 4756 3187
rect 4722 3059 4756 3099
rect 4722 2979 4756 3019
rect 4722 2899 4756 2939
rect 4722 2819 4756 2859
rect 3252 2660 3286 2700
rect 3252 2580 3286 2620
rect 3252 2500 3286 2540
rect 3252 2420 3286 2460
rect 3252 2340 3286 2380
rect 4722 2739 4756 2779
rect 4722 2659 4756 2699
rect 4722 2579 4756 2619
rect 4722 2499 4756 2539
rect 4722 2411 4756 2459
rect 5140 3139 5174 3187
rect 5140 3059 5174 3099
rect 5140 2979 5174 3019
rect 5140 2899 5174 2939
rect 5140 2819 5174 2859
rect 5140 2739 5174 2779
rect 5140 2659 5174 2699
rect 5140 2579 5174 2619
rect 5140 2499 5174 2539
rect 5140 2411 5174 2459
rect 5558 3139 5592 3187
rect 5558 3059 5592 3099
rect 5558 2979 5592 3019
rect 5558 2899 5592 2939
rect 5558 2819 5592 2859
rect 5558 2739 5592 2779
rect 5558 2659 5592 2699
rect 5558 2579 5592 2619
rect 5558 2499 5592 2539
rect 5558 2411 5592 2459
rect 250 982 284 1022
rect 250 902 284 942
rect 250 822 284 862
rect 250 742 284 782
rect 250 662 284 702
rect 250 582 284 622
rect 250 502 284 542
rect 250 422 284 462
rect 250 342 284 382
rect 250 262 284 302
rect 250 172 284 222
rect 668 970 702 1010
rect 668 890 702 930
rect 668 810 702 850
rect 668 730 702 770
rect 668 650 702 690
rect 668 570 702 610
rect 668 490 702 530
rect 668 410 702 450
rect 668 330 702 370
rect 668 250 702 290
rect 668 172 702 210
rect 1086 982 1120 1022
rect 1086 902 1120 942
rect 1086 822 1120 862
rect 1086 742 1120 782
rect 1086 662 1120 702
rect 1086 582 1120 622
rect 1086 502 1120 542
rect 1086 422 1120 462
rect 1086 342 1120 382
rect 1086 262 1120 302
rect 1086 172 1120 222
rect 1504 982 1538 1048
rect 1504 902 1538 942
rect 1504 822 1538 862
rect 1504 742 1538 782
rect 1504 662 1538 702
rect 1504 582 1538 622
rect 1504 502 1538 542
rect 1504 422 1538 462
rect 1504 342 1538 382
rect 1504 262 1538 302
rect 1504 172 1538 222
rect 1922 982 1956 1048
rect 1922 902 1956 942
rect 1922 822 1956 862
rect 1922 742 1956 782
rect 1922 662 1956 702
rect 1922 582 1956 622
rect 3845 902 3879 950
rect 3845 822 3879 862
rect 3845 742 3879 782
rect 3845 662 3879 702
rect 3845 582 3879 622
rect 1922 502 1956 542
rect 1922 422 1956 462
rect 1922 342 1956 382
rect 1922 262 1956 302
rect 1922 172 1956 222
rect 3845 502 3879 542
rect 3845 422 3879 462
rect 3845 342 3879 382
rect 3845 262 3879 302
rect 3845 174 3879 222
rect 4263 902 4297 950
rect 4263 822 4297 862
rect 4263 742 4297 782
rect 4263 662 4297 702
rect 4263 582 4297 622
rect 4263 502 4297 542
rect 4263 422 4297 462
rect 4263 342 4297 382
rect 4263 262 4297 302
rect 4263 174 4297 222
rect 4681 902 4715 950
rect 4681 822 4715 862
rect 4681 742 4715 782
rect 4681 662 4715 702
rect 4681 582 4715 622
rect 4681 502 4715 542
rect 4681 422 4715 462
rect 4681 342 4715 382
rect 4681 262 4715 302
rect 4681 174 4715 222
<< pdiffc >>
rect 250 2600 284 2642
rect 250 2520 284 2560
rect 250 2440 284 2480
rect 250 2360 284 2400
rect 250 2280 284 2320
rect 250 2200 284 2240
rect 250 2120 284 2160
rect 250 2040 284 2080
rect 250 1960 284 2000
rect 250 1880 284 1920
rect 250 1800 284 1840
rect 668 2568 702 2608
rect 668 2488 702 2528
rect 668 2408 702 2448
rect 668 2328 702 2368
rect 668 2248 702 2288
rect 668 2168 702 2208
rect 668 2088 702 2128
rect 668 2008 702 2048
rect 668 1928 702 1968
rect 668 1848 702 1888
rect 668 1766 702 1808
rect 1086 2600 1120 2642
rect 1086 2520 1120 2560
rect 1086 2440 1120 2480
rect 1086 2360 1120 2400
rect 1086 2280 1120 2320
rect 1086 2200 1120 2240
rect 1086 2120 1120 2160
rect 1086 2040 1120 2080
rect 1086 1960 1120 2000
rect 1086 1880 1120 1920
rect 1086 1800 1120 1840
rect 3845 2580 3879 2631
rect 3845 2500 3879 2540
rect 3845 2420 3879 2460
rect 3845 2340 3879 2380
rect 3845 2260 3879 2300
rect 3845 2180 3879 2220
rect 3845 2100 3879 2140
rect 3845 2020 3879 2060
rect 3845 1922 3879 1980
rect 4263 2580 4297 2631
rect 4263 2500 4297 2540
rect 4263 2420 4297 2460
rect 4263 2340 4297 2380
rect 4263 2260 4297 2300
rect 4263 2180 4297 2220
rect 4263 2100 4297 2140
rect 4263 2020 4297 2060
rect 4263 1940 4297 1980
rect 4263 1855 4297 1900
rect 2416 1512 2450 1552
rect 2416 1432 2450 1472
rect 2416 1352 2450 1392
rect 2416 1272 2450 1312
rect 2416 1192 2450 1232
rect 2416 1112 2450 1152
rect 2416 1032 2450 1072
rect 2416 952 2450 992
rect 2416 872 2450 912
rect 2416 792 2450 832
rect 2416 710 2450 752
rect 2834 1544 2868 1586
rect 2834 1464 2868 1504
rect 2834 1384 2868 1424
rect 2834 1304 2868 1344
rect 2834 1224 2868 1264
rect 2834 1144 2868 1184
rect 2834 1064 2868 1104
rect 2834 984 2868 1024
rect 2834 904 2868 944
rect 2834 824 2868 864
rect 2834 744 2868 784
rect 3252 1512 3286 1552
rect 3252 1432 3286 1472
rect 3252 1352 3286 1392
rect 3252 1272 3286 1312
rect 3252 1192 3286 1232
rect 3252 1112 3286 1152
rect 3252 1032 3286 1072
rect 3252 952 3286 992
rect 3252 872 3286 912
rect 3252 792 3286 832
rect 3252 710 3286 752
rect 5140 1462 5174 1506
rect 5140 1382 5174 1422
rect 5140 1302 5174 1342
rect 5140 1222 5174 1262
rect 5140 1142 5174 1182
rect 5140 1062 5174 1102
rect 5140 982 5174 1022
rect 5140 902 5174 942
rect 5140 822 5174 862
rect 5140 730 5174 782
rect 5558 1462 5592 1506
rect 5558 1382 5592 1422
rect 5558 1302 5592 1342
rect 5558 1222 5592 1262
rect 5558 1142 5592 1182
rect 5558 1062 5592 1102
rect 5558 982 5592 1022
rect 5558 902 5592 942
rect 5558 822 5592 862
rect 5558 730 5592 782
<< nsubdiff >>
rect 136 2745 232 2779
rect 280 2745 320 2779
rect 360 2745 400 2779
rect 440 2745 480 2779
rect 520 2745 560 2779
rect 600 2745 640 2779
rect 680 2745 720 2779
rect 760 2745 800 2779
rect 840 2745 880 2779
rect 920 2745 960 2779
rect 1000 2745 1040 2779
rect 1100 2745 1234 2779
rect 136 2693 170 2745
rect 1200 2694 1234 2745
rect 136 2600 170 2640
rect 136 2520 170 2560
rect 136 2440 170 2480
rect 136 2360 170 2400
rect 136 2280 170 2320
rect 136 2200 170 2240
rect 136 2120 170 2160
rect 136 2040 170 2080
rect 136 1960 170 2000
rect 136 1880 170 1920
rect 136 1749 170 1820
rect 1200 2620 1234 2660
rect 1200 2540 1234 2580
rect 1200 2460 1234 2500
rect 1200 2380 1234 2420
rect 1200 2300 1234 2340
rect 3731 2744 3827 2778
rect 3880 2744 3920 2778
rect 3960 2744 4000 2778
rect 4040 2744 4080 2778
rect 4120 2744 4160 2778
rect 4200 2744 4240 2778
rect 4315 2744 4411 2778
rect 3731 2730 3765 2744
rect 4377 2730 4411 2744
rect 3731 2638 3765 2678
rect 3731 2558 3765 2598
rect 3731 2478 3765 2518
rect 3731 2398 3765 2438
rect 3731 2318 3765 2358
rect 1200 2220 1234 2260
rect 1200 2140 1234 2180
rect 1200 2060 1234 2100
rect 1200 1980 1234 2020
rect 1200 1900 1234 1940
rect 1200 1820 1234 1860
rect 1200 1749 1234 1785
rect 3731 2238 3765 2278
rect 3731 2158 3765 2198
rect 3731 2078 3765 2118
rect 3731 1998 3765 2038
rect 3731 1935 3765 1964
rect 4377 2640 4411 2680
rect 4377 2560 4411 2600
rect 4377 2480 4411 2520
rect 4377 2400 4411 2440
rect 4377 2320 4411 2360
rect 4377 2240 4411 2280
rect 4377 2160 4411 2200
rect 4377 2080 4411 2120
rect 4377 2000 4411 2040
rect 4377 1937 4411 1966
rect 2302 1533 2336 1572
rect 2302 1458 2336 1498
rect 2302 1378 2336 1418
rect 2302 1298 2336 1338
rect 2302 1218 2336 1258
rect 2302 1138 2336 1178
rect 2302 1058 2336 1098
rect 2302 978 2336 1018
rect 2302 898 2336 938
rect 2302 818 2336 858
rect 2302 738 2336 778
rect 3366 1532 3400 1560
rect 3366 1432 3400 1472
rect 3366 1352 3400 1392
rect 3366 1272 3400 1312
rect 3366 1192 3400 1232
rect 3366 1112 3400 1152
rect 3366 1032 3400 1072
rect 3366 952 3400 992
rect 5026 1172 5060 1212
rect 5026 1092 5060 1132
rect 5026 1012 5060 1052
rect 3366 872 3400 912
rect 3366 792 3400 832
rect 3366 712 3400 752
rect 2302 658 2336 698
rect 2302 607 2336 624
rect 3366 607 3400 659
rect 2302 573 2436 607
rect 2496 573 2536 607
rect 2576 573 2616 607
rect 2656 573 2696 607
rect 2736 573 2776 607
rect 2816 573 2856 607
rect 2896 573 2936 607
rect 2976 573 3016 607
rect 3056 573 3096 607
rect 3136 573 3176 607
rect 3216 573 3256 607
rect 3304 573 3400 607
rect 5026 932 5060 972
rect 5026 852 5060 892
rect 5026 772 5060 812
rect 5026 692 5060 732
rect 5672 1493 5706 1523
rect 5672 1410 5706 1450
rect 5672 1330 5706 1370
rect 5672 1250 5706 1290
rect 5672 1170 5706 1210
rect 5672 1090 5706 1130
rect 5672 1010 5706 1050
rect 5672 930 5706 970
rect 5672 850 5706 890
rect 5672 770 5706 810
rect 5672 690 5706 730
rect 5026 583 5060 652
rect 5672 617 5706 631
rect 5120 583 5160 617
rect 5200 583 5240 617
rect 5280 583 5320 617
rect 5360 583 5400 617
rect 5440 583 5480 617
rect 5520 583 5560 617
rect 5610 583 5706 617
<< nsubdiffcont >>
rect 232 2745 280 2779
rect 320 2745 360 2779
rect 400 2745 440 2779
rect 480 2745 520 2779
rect 560 2745 600 2779
rect 640 2745 680 2779
rect 720 2745 760 2779
rect 800 2745 840 2779
rect 880 2745 920 2779
rect 960 2745 1000 2779
rect 1040 2745 1100 2779
rect 136 2640 170 2693
rect 1200 2660 1234 2694
rect 136 2560 170 2600
rect 136 2480 170 2520
rect 136 2400 170 2440
rect 136 2320 170 2360
rect 136 2240 170 2280
rect 136 2160 170 2200
rect 136 2080 170 2120
rect 136 2000 170 2040
rect 136 1920 170 1960
rect 136 1820 170 1880
rect 1200 2580 1234 2620
rect 1200 2500 1234 2540
rect 1200 2420 1234 2460
rect 1200 2340 1234 2380
rect 3827 2744 3880 2778
rect 3920 2744 3960 2778
rect 4000 2744 4040 2778
rect 4080 2744 4120 2778
rect 4160 2744 4200 2778
rect 4240 2744 4315 2778
rect 3731 2678 3765 2730
rect 4377 2680 4411 2730
rect 3731 2598 3765 2638
rect 3731 2518 3765 2558
rect 3731 2438 3765 2478
rect 3731 2358 3765 2398
rect 1200 2260 1234 2300
rect 1200 2180 1234 2220
rect 1200 2100 1234 2140
rect 1200 2020 1234 2060
rect 1200 1940 1234 1980
rect 1200 1860 1234 1900
rect 1200 1785 1234 1820
rect 3731 2278 3765 2318
rect 3731 2198 3765 2238
rect 3731 2118 3765 2158
rect 3731 2038 3765 2078
rect 3731 1964 3765 1998
rect 4377 2600 4411 2640
rect 4377 2520 4411 2560
rect 4377 2440 4411 2480
rect 4377 2360 4411 2400
rect 4377 2280 4411 2320
rect 4377 2200 4411 2240
rect 4377 2120 4411 2160
rect 4377 2040 4411 2080
rect 4377 1966 4411 2000
rect 2302 1498 2336 1533
rect 2302 1418 2336 1458
rect 2302 1338 2336 1378
rect 2302 1258 2336 1298
rect 2302 1178 2336 1218
rect 2302 1098 2336 1138
rect 2302 1018 2336 1058
rect 2302 938 2336 978
rect 2302 858 2336 898
rect 2302 778 2336 818
rect 2302 698 2336 738
rect 3366 1472 3400 1532
rect 3366 1392 3400 1432
rect 3366 1312 3400 1352
rect 3366 1232 3400 1272
rect 3366 1152 3400 1192
rect 3366 1072 3400 1112
rect 3366 992 3400 1032
rect 5026 1132 5060 1172
rect 5026 1052 5060 1092
rect 5026 972 5060 1012
rect 3366 912 3400 952
rect 3366 832 3400 872
rect 3366 752 3400 792
rect 2302 624 2336 658
rect 3366 659 3400 712
rect 2436 573 2496 607
rect 2536 573 2576 607
rect 2616 573 2656 607
rect 2696 573 2736 607
rect 2776 573 2816 607
rect 2856 573 2896 607
rect 2936 573 2976 607
rect 3016 573 3056 607
rect 3096 573 3136 607
rect 3176 573 3216 607
rect 3256 573 3304 607
rect 5026 892 5060 932
rect 5026 812 5060 852
rect 5026 732 5060 772
rect 5672 1450 5706 1493
rect 5672 1370 5706 1410
rect 5672 1290 5706 1330
rect 5672 1210 5706 1250
rect 5672 1130 5706 1170
rect 5672 1050 5706 1090
rect 5672 970 5706 1010
rect 5672 890 5706 930
rect 5672 810 5706 850
rect 5672 730 5706 770
rect 5026 652 5060 692
rect 5672 631 5706 690
rect 5060 583 5120 617
rect 5160 583 5200 617
rect 5240 583 5280 617
rect 5320 583 5360 617
rect 5400 583 5440 617
rect 5480 583 5520 617
rect 5560 583 5610 617
<< poly >>
rect 1626 3202 1986 3242
rect 2044 3202 2404 3242
rect 2462 3202 2822 3242
rect 2880 3202 3240 3242
rect 296 2654 656 2680
rect 714 2654 1074 2680
rect 4768 3199 5128 3239
rect 5186 3199 5546 3239
rect 3891 2643 4251 2683
rect 1626 2214 1986 2302
rect 2044 2214 2404 2302
rect 2462 2214 2822 2302
rect 2880 2214 3240 2302
rect 1626 2140 3240 2214
rect 1626 2088 3020 2140
rect 296 1692 656 1754
rect 714 1692 1074 1754
rect 2600 2040 3020 2088
rect 3100 2040 3140 2140
rect 3220 2040 3240 2140
rect 2600 2000 3240 2040
rect 2600 1880 2616 2000
rect 2736 1880 2776 2000
rect 2896 1880 2936 2000
rect 3056 1880 3096 2000
rect 3216 1880 3240 2000
rect 2600 1748 3240 1880
rect 4768 2339 5128 2399
rect 5186 2339 5546 2399
rect 4768 2139 5546 2339
rect 5185 2060 5546 2139
rect 5185 1972 5326 2060
rect 5406 1972 5446 2060
rect 5526 1972 5546 2060
rect 5185 1938 5546 1972
rect 5185 1858 5326 1938
rect 5406 1858 5446 1938
rect 5526 1858 5546 1938
rect 296 1552 1074 1692
rect 2462 1664 3240 1748
rect 2462 1598 2822 1664
rect 2880 1598 3240 1664
rect 296 1516 936 1552
rect 286 1506 936 1516
rect 286 1426 296 1506
rect 376 1426 410 1506
rect 490 1426 936 1506
rect 286 1390 936 1426
rect 286 1306 296 1390
rect 376 1306 410 1390
rect 490 1314 936 1390
rect 490 1306 1910 1314
rect 286 1296 1910 1306
rect 296 1148 1910 1296
rect 296 1060 656 1148
rect 714 1060 1074 1148
rect 1132 1060 1492 1148
rect 1550 1060 1910 1148
rect 3891 1496 4251 1843
rect 5185 1615 5546 1858
rect 5186 1518 5546 1615
rect 3891 1416 3902 1496
rect 3982 1416 4028 1496
rect 4108 1416 4251 1496
rect 3891 1382 4251 1416
rect 3891 1302 3902 1382
rect 3982 1302 4028 1382
rect 4108 1302 4251 1382
rect 3891 1222 4251 1302
rect 3891 1022 4669 1222
rect 3891 962 4251 1022
rect 4309 962 4669 1022
rect 2462 672 2822 698
rect 2880 672 3240 698
rect 5186 678 5546 718
rect 296 120 656 160
rect 714 120 1074 160
rect 1132 120 1492 160
rect 1550 120 1910 160
rect 3891 122 4251 162
rect 4309 122 4669 162
<< polycont >>
rect 3020 2040 3100 2140
rect 3140 2040 3220 2140
rect 2616 1880 2736 2000
rect 2776 1880 2896 2000
rect 2936 1880 3056 2000
rect 3096 1880 3216 2000
rect 5326 1972 5406 2060
rect 5446 1972 5526 2060
rect 5326 1858 5406 1938
rect 5446 1858 5526 1938
rect 296 1426 376 1506
rect 410 1426 490 1506
rect 296 1306 376 1390
rect 410 1306 490 1390
rect 3902 1416 3982 1496
rect 4028 1416 4108 1496
rect 3902 1302 3982 1382
rect 4028 1302 4108 1382
<< locali >>
rect 1466 3354 1936 3360
rect 1569 3270 1607 3354
rect 1691 3270 1729 3354
rect 1813 3270 1851 3354
rect 1935 3270 1936 3354
rect 1466 3264 1936 3270
rect 2146 3354 2718 3360
rect 2230 3270 2268 3354
rect 2352 3270 2390 3354
rect 2474 3270 2512 3354
rect 2596 3270 2634 3354
rect 2146 3264 2718 3270
rect 2931 3354 3400 3360
rect 3015 3270 3053 3354
rect 3137 3270 3175 3354
rect 3259 3270 3297 3354
rect 2931 3264 3400 3270
rect 4608 3354 5076 3360
rect 5238 3354 5706 3360
rect 4710 3270 4750 3354
rect 4832 3270 4872 3354
rect 4954 3270 4994 3354
rect 5321 3270 5359 3354
rect 5443 3270 5481 3354
rect 5565 3270 5603 3354
rect 4608 3264 5076 3270
rect 5238 3264 5706 3270
rect 1568 3190 1626 3264
rect 1568 3140 1580 3190
rect 1614 3140 1626 3190
rect 1568 3100 1626 3140
rect 1568 3060 1580 3100
rect 1614 3060 1626 3100
rect 1568 3020 1626 3060
rect 1568 2980 1580 3020
rect 1614 2980 1626 3020
rect 1568 2940 1626 2980
rect 1568 2900 1580 2940
rect 1614 2900 1626 2940
rect 1568 2860 1626 2900
rect 1568 2820 1580 2860
rect 1614 2820 1626 2860
rect 136 2810 605 2816
rect 239 2779 277 2810
rect 239 2726 277 2745
rect 361 2726 399 2810
rect 483 2779 521 2810
rect 765 2810 1234 2816
rect 765 2779 801 2810
rect 885 2779 923 2810
rect 1007 2779 1045 2810
rect 520 2745 521 2779
rect 605 2745 640 2779
rect 680 2745 720 2779
rect 760 2745 800 2779
rect 920 2745 923 2779
rect 1007 2745 1040 2779
rect 483 2726 521 2745
rect 136 2720 605 2726
rect 765 2726 801 2745
rect 885 2726 923 2745
rect 1007 2726 1045 2745
rect 1129 2726 1167 2810
rect 1568 2780 1626 2820
rect 1568 2740 1580 2780
rect 1614 2740 1626 2780
rect 765 2720 1234 2726
rect 136 2693 170 2720
rect 136 2600 170 2640
rect 136 2520 170 2560
rect 136 2440 170 2480
rect 136 2360 170 2400
rect 136 2280 170 2320
rect 136 2200 170 2240
rect 136 2120 170 2160
rect 136 2040 170 2080
rect 136 1960 170 2000
rect 136 1880 170 1920
rect 136 1749 170 1820
rect 238 2642 296 2720
rect 238 2600 250 2642
rect 284 2600 296 2642
rect 238 2560 296 2600
rect 238 2520 250 2560
rect 284 2520 296 2560
rect 238 2480 296 2520
rect 238 2440 250 2480
rect 284 2440 296 2480
rect 238 2400 296 2440
rect 238 2360 250 2400
rect 284 2360 296 2400
rect 238 2320 296 2360
rect 238 2280 250 2320
rect 284 2280 296 2320
rect 238 2240 296 2280
rect 238 2200 250 2240
rect 284 2200 296 2240
rect 238 2160 296 2200
rect 238 2120 250 2160
rect 284 2120 296 2160
rect 238 2080 296 2120
rect 238 2040 250 2080
rect 284 2040 296 2080
rect 238 2000 296 2040
rect 238 1960 250 2000
rect 284 1960 296 2000
rect 238 1920 296 1960
rect 238 1880 250 1920
rect 284 1880 296 1920
rect 238 1840 296 1880
rect 238 1800 250 1840
rect 284 1800 296 1840
rect 238 1750 296 1800
rect 656 2608 714 2658
rect 656 2568 668 2608
rect 702 2568 714 2608
rect 656 2528 714 2568
rect 656 2488 668 2528
rect 702 2488 714 2528
rect 656 2448 714 2488
rect 656 2408 668 2448
rect 702 2408 714 2448
rect 656 2368 714 2408
rect 656 2328 668 2368
rect 702 2328 714 2368
rect 656 2288 714 2328
rect 656 2248 668 2288
rect 702 2248 714 2288
rect 656 2208 714 2248
rect 656 2168 668 2208
rect 702 2168 714 2208
rect 656 2128 714 2168
rect 656 2088 668 2128
rect 702 2088 714 2128
rect 656 2048 714 2088
rect 656 2008 668 2048
rect 702 2008 714 2048
rect 656 1968 714 2008
rect 656 1928 668 1968
rect 702 1928 714 1968
rect 656 1888 714 1928
rect 656 1848 668 1888
rect 702 1848 714 1888
rect 656 1808 714 1848
rect 656 1766 668 1808
rect 702 1766 714 1808
rect 280 1500 296 1506
rect 376 1500 410 1506
rect 280 1312 286 1500
rect 490 1426 506 1506
rect 488 1390 506 1426
rect 280 1306 296 1312
rect 376 1306 410 1312
rect 490 1306 506 1390
rect 656 1468 714 1766
rect 1074 2642 1132 2720
rect 1074 2600 1086 2642
rect 1120 2600 1132 2642
rect 1074 2560 1132 2600
rect 1074 2520 1086 2560
rect 1120 2520 1132 2560
rect 1074 2480 1132 2520
rect 1074 2440 1086 2480
rect 1120 2440 1132 2480
rect 1074 2400 1132 2440
rect 1074 2360 1086 2400
rect 1120 2360 1132 2400
rect 1074 2320 1132 2360
rect 1074 2280 1086 2320
rect 1120 2280 1132 2320
rect 1074 2240 1132 2280
rect 1074 2200 1086 2240
rect 1120 2200 1132 2240
rect 1074 2160 1132 2200
rect 1074 2120 1086 2160
rect 1120 2120 1132 2160
rect 1074 2080 1132 2120
rect 1074 2040 1086 2080
rect 1120 2040 1132 2080
rect 1074 2000 1132 2040
rect 1074 1960 1086 2000
rect 1120 1960 1132 2000
rect 1074 1920 1132 1960
rect 1074 1880 1086 1920
rect 1120 1880 1132 1920
rect 1074 1840 1132 1880
rect 1074 1800 1086 1840
rect 1120 1800 1132 1840
rect 1074 1750 1132 1800
rect 1200 2694 1234 2720
rect 1200 2620 1234 2660
rect 1200 2540 1234 2580
rect 1200 2460 1234 2500
rect 1200 2380 1234 2420
rect 1568 2700 1626 2740
rect 1568 2660 1580 2700
rect 1614 2660 1626 2700
rect 1568 2620 1626 2660
rect 1568 2580 1580 2620
rect 1614 2580 1626 2620
rect 1568 2540 1626 2580
rect 1568 2500 1580 2540
rect 1614 2500 1626 2540
rect 1568 2460 1626 2500
rect 1568 2420 1580 2460
rect 1614 2420 1626 2460
rect 1568 2380 1626 2420
rect 1568 2347 1580 2380
rect 1575 2345 1580 2347
rect 1200 2300 1234 2340
rect 1614 2347 1626 2380
rect 1986 3190 2044 3206
rect 1986 3140 1998 3190
rect 2032 3140 2044 3190
rect 1986 3100 2044 3140
rect 1986 3060 1998 3100
rect 2032 3060 2044 3100
rect 1986 3020 2044 3060
rect 1986 2980 1998 3020
rect 2032 2980 2044 3020
rect 1986 2940 2044 2980
rect 1986 2900 1998 2940
rect 2032 2900 2044 2940
rect 1986 2860 2044 2900
rect 1986 2820 1998 2860
rect 2032 2820 2044 2860
rect 1986 2780 2044 2820
rect 1986 2740 1998 2780
rect 2032 2740 2044 2780
rect 1986 2700 2044 2740
rect 1986 2660 1998 2700
rect 2032 2660 2044 2700
rect 1986 2620 2044 2660
rect 1986 2580 1998 2620
rect 2032 2580 2044 2620
rect 1986 2540 2044 2580
rect 1986 2500 1998 2540
rect 2032 2500 2044 2540
rect 1986 2460 2044 2500
rect 1986 2420 1998 2460
rect 2032 2420 2044 2460
rect 1986 2380 2044 2420
rect 1580 2298 1614 2314
rect 1986 2314 1998 2380
rect 2032 2314 2044 2380
rect 2404 3190 2462 3264
rect 2404 3140 2416 3190
rect 2450 3140 2462 3190
rect 2404 3100 2462 3140
rect 2404 3060 2416 3100
rect 2450 3060 2462 3100
rect 2404 3020 2462 3060
rect 2404 2980 2416 3020
rect 2450 2980 2462 3020
rect 2404 2940 2462 2980
rect 2404 2900 2416 2940
rect 2450 2900 2462 2940
rect 2404 2860 2462 2900
rect 2404 2820 2416 2860
rect 2450 2820 2462 2860
rect 2404 2780 2462 2820
rect 2404 2740 2416 2780
rect 2450 2740 2462 2780
rect 2404 2700 2462 2740
rect 2404 2660 2416 2700
rect 2450 2660 2462 2700
rect 2404 2620 2462 2660
rect 2404 2580 2416 2620
rect 2450 2580 2462 2620
rect 2404 2540 2462 2580
rect 2404 2500 2416 2540
rect 2450 2500 2462 2540
rect 2404 2460 2462 2500
rect 2404 2420 2416 2460
rect 2450 2420 2462 2460
rect 2404 2380 2462 2420
rect 2404 2347 2416 2380
rect 1200 2220 1234 2260
rect 1200 2140 1234 2180
rect 1200 2060 1234 2100
rect 1986 2140 2044 2314
rect 2450 2347 2462 2380
rect 2822 3190 2880 3206
rect 2822 3152 2834 3190
rect 2868 3152 2880 3190
rect 2822 3112 2880 3152
rect 2822 3072 2834 3112
rect 2868 3072 2880 3112
rect 2822 3032 2880 3072
rect 2822 2992 2834 3032
rect 2868 2992 2880 3032
rect 2822 2952 2880 2992
rect 2822 2912 2834 2952
rect 2868 2912 2880 2952
rect 2822 2872 2880 2912
rect 2822 2832 2834 2872
rect 2868 2832 2880 2872
rect 2822 2792 2880 2832
rect 2822 2752 2834 2792
rect 2868 2752 2880 2792
rect 2822 2712 2880 2752
rect 2822 2672 2834 2712
rect 2868 2672 2880 2712
rect 2822 2632 2880 2672
rect 2822 2592 2834 2632
rect 2868 2592 2880 2632
rect 2822 2552 2880 2592
rect 2822 2512 2834 2552
rect 2868 2512 2880 2552
rect 2822 2472 2880 2512
rect 2822 2432 2834 2472
rect 2868 2432 2880 2472
rect 2822 2392 2880 2432
rect 2822 2352 2834 2392
rect 2868 2352 2880 2392
rect 2416 2302 2450 2340
rect 2822 2140 2880 2352
rect 3240 3190 3298 3264
rect 3240 3140 3252 3190
rect 3286 3140 3298 3190
rect 3240 3100 3298 3140
rect 3240 3060 3252 3100
rect 3286 3060 3298 3100
rect 3240 3020 3298 3060
rect 3240 2980 3252 3020
rect 3286 2980 3298 3020
rect 3240 2940 3298 2980
rect 3240 2900 3252 2940
rect 3286 2900 3298 2940
rect 3240 2860 3298 2900
rect 3240 2820 3252 2860
rect 3286 2820 3298 2860
rect 3240 2780 3298 2820
rect 4710 3187 4768 3264
rect 4710 3139 4722 3187
rect 4756 3139 4768 3187
rect 4710 3099 4768 3139
rect 4710 3059 4722 3099
rect 4756 3059 4768 3099
rect 4710 3019 4768 3059
rect 4710 2979 4722 3019
rect 4756 2979 4768 3019
rect 4710 2939 4768 2979
rect 4710 2899 4722 2939
rect 4756 2899 4768 2939
rect 4710 2859 4768 2899
rect 4710 2819 4722 2859
rect 4756 2819 4768 2859
rect 3240 2740 3252 2780
rect 3286 2740 3298 2780
rect 3240 2700 3298 2740
rect 3240 2660 3252 2700
rect 3286 2660 3298 2700
rect 3240 2620 3298 2660
rect 3240 2580 3252 2620
rect 3286 2580 3298 2620
rect 3240 2540 3298 2580
rect 3240 2500 3252 2540
rect 3286 2500 3298 2540
rect 3240 2460 3298 2500
rect 3240 2420 3252 2460
rect 3286 2420 3298 2460
rect 3240 2380 3298 2420
rect 3240 2347 3252 2380
rect 3286 2347 3298 2380
rect 3731 2810 4150 2816
rect 3815 2778 3853 2810
rect 3937 2778 3975 2810
rect 4059 2778 4097 2810
rect 4710 2779 4768 2819
rect 3815 2744 3827 2778
rect 3960 2744 3975 2778
rect 4059 2744 4080 2778
rect 4200 2744 4240 2778
rect 4315 2744 4411 2778
rect 3815 2726 3853 2744
rect 3937 2726 3975 2744
rect 4059 2726 4097 2744
rect 4377 2730 4411 2744
rect 3765 2720 4150 2726
rect 3731 2638 3765 2678
rect 3731 2558 3765 2598
rect 3731 2478 3765 2518
rect 3731 2398 3765 2438
rect 3252 2302 3286 2340
rect 3731 2318 3765 2358
rect 3731 2238 3765 2278
rect 3731 2158 3765 2198
rect 1986 2082 2880 2140
rect 1200 1980 1234 2020
rect 1200 1900 1234 1940
rect 1200 1820 1234 1860
rect 1200 1749 1234 1785
rect 2294 1794 2394 2082
rect 3000 2040 3020 2140
rect 3100 2040 3140 2140
rect 3220 2040 3240 2140
rect 3000 2024 3240 2040
rect 3731 2078 3765 2118
rect 3000 2018 3400 2024
rect 3000 2000 3080 2018
rect 2736 1880 2760 2000
rect 2896 1880 2920 2000
rect 3056 1880 3080 2000
rect 3220 1892 3260 2018
rect 3388 1892 3400 2018
rect 3731 1998 3765 2038
rect 3731 1935 3765 1964
rect 3833 2631 3891 2720
rect 3833 2580 3845 2631
rect 3879 2580 3891 2631
rect 3833 2540 3891 2580
rect 3833 2500 3845 2540
rect 3879 2500 3891 2540
rect 3833 2460 3891 2500
rect 3833 2420 3845 2460
rect 3879 2420 3891 2460
rect 3833 2380 3891 2420
rect 3833 2340 3845 2380
rect 3879 2340 3891 2380
rect 3833 2300 3891 2340
rect 3833 2260 3845 2300
rect 3879 2260 3891 2300
rect 3833 2220 3891 2260
rect 3833 2180 3845 2220
rect 3879 2180 3891 2220
rect 3833 2140 3891 2180
rect 3833 2100 3845 2140
rect 3879 2100 3891 2140
rect 3833 2060 3891 2100
rect 3833 2020 3845 2060
rect 3879 2020 3891 2060
rect 3833 1980 3891 2020
rect 3833 1922 3845 1980
rect 3879 1922 3891 1980
rect 3833 1906 3891 1922
rect 4251 2631 4310 2647
rect 4251 2580 4263 2631
rect 4297 2580 4310 2631
rect 4251 2540 4310 2580
rect 4251 2500 4263 2540
rect 4297 2500 4310 2540
rect 4251 2460 4310 2500
rect 4251 2420 4263 2460
rect 4297 2420 4310 2460
rect 4251 2380 4310 2420
rect 4251 2340 4263 2380
rect 4297 2340 4310 2380
rect 4251 2300 4310 2340
rect 4251 2260 4263 2300
rect 4297 2260 4310 2300
rect 4251 2220 4310 2260
rect 4251 2180 4263 2220
rect 4297 2180 4310 2220
rect 4251 2140 4310 2180
rect 4251 2100 4263 2140
rect 4297 2100 4310 2140
rect 4251 2060 4310 2100
rect 4251 2020 4263 2060
rect 4297 2020 4310 2060
rect 4251 1980 4310 2020
rect 4251 1940 4263 1980
rect 4297 1940 4310 1980
rect 3220 1880 3400 1892
rect 4251 1900 4310 1940
rect 4377 2640 4411 2680
rect 4377 2560 4411 2600
rect 4377 2480 4411 2520
rect 4377 2400 4411 2440
rect 4710 2739 4722 2779
rect 4756 2739 4768 2779
rect 4710 2699 4768 2739
rect 4710 2659 4722 2699
rect 4756 2659 4768 2699
rect 4710 2619 4768 2659
rect 4710 2579 4722 2619
rect 4756 2579 4768 2619
rect 4710 2539 4768 2579
rect 4710 2499 4722 2539
rect 4756 2499 4768 2539
rect 4710 2459 4768 2499
rect 4710 2411 4722 2459
rect 4756 2411 4768 2459
rect 4710 2395 4768 2411
rect 5127 3187 5186 3203
rect 5127 3139 5140 3187
rect 5174 3139 5186 3187
rect 5127 3099 5186 3139
rect 5127 3059 5140 3099
rect 5174 3059 5186 3099
rect 5127 3019 5186 3059
rect 5127 2979 5140 3019
rect 5174 2979 5186 3019
rect 5127 2939 5186 2979
rect 5127 2899 5140 2939
rect 5174 2899 5186 2939
rect 5127 2859 5186 2899
rect 5127 2819 5140 2859
rect 5174 2819 5186 2859
rect 5127 2779 5186 2819
rect 5127 2739 5140 2779
rect 5174 2739 5186 2779
rect 5127 2699 5186 2739
rect 5127 2659 5140 2699
rect 5174 2659 5186 2699
rect 5127 2619 5186 2659
rect 5127 2579 5140 2619
rect 5174 2579 5186 2619
rect 5127 2539 5186 2579
rect 5127 2499 5140 2539
rect 5174 2499 5186 2539
rect 5127 2459 5186 2499
rect 5127 2411 5140 2459
rect 5174 2411 5186 2459
rect 4377 2320 4411 2360
rect 4377 2240 4411 2280
rect 4377 2160 4411 2200
rect 4377 2080 4411 2120
rect 4377 2000 4411 2040
rect 4377 1937 4411 1966
rect 4713 2012 4813 2024
rect 4251 1855 4263 1900
rect 4297 1855 4310 1900
rect 4251 1794 4310 1855
rect 4713 1794 4813 1892
rect 2294 1694 4813 1794
rect 2302 1533 2336 1572
rect 656 1368 1492 1468
rect 250 1022 284 1064
rect 238 982 250 1015
rect 284 982 296 1015
rect 238 942 296 982
rect 238 902 250 942
rect 284 902 296 942
rect 238 862 296 902
rect 238 822 250 862
rect 284 822 296 862
rect 238 782 296 822
rect 238 742 250 782
rect 284 742 296 782
rect 238 702 296 742
rect 238 662 250 702
rect 284 662 296 702
rect 238 622 296 662
rect 238 582 250 622
rect 284 582 296 622
rect 238 542 296 582
rect 238 502 250 542
rect 284 502 296 542
rect 238 462 296 502
rect 238 422 250 462
rect 284 422 296 462
rect 238 382 296 422
rect 238 342 250 382
rect 284 342 296 382
rect 238 302 296 342
rect 238 262 250 302
rect 284 262 296 302
rect 238 222 296 262
rect 238 172 250 222
rect 284 172 296 222
rect 238 96 296 172
rect 656 1010 714 1368
rect 2302 1458 2336 1498
rect 2302 1378 2336 1418
rect 1086 1022 1120 1064
rect 656 970 668 1010
rect 702 970 714 1010
rect 656 930 714 970
rect 656 890 668 930
rect 702 890 714 930
rect 656 850 714 890
rect 656 810 668 850
rect 702 810 714 850
rect 656 770 714 810
rect 656 730 668 770
rect 702 730 714 770
rect 656 690 714 730
rect 656 650 668 690
rect 702 650 714 690
rect 656 610 714 650
rect 656 570 668 610
rect 702 570 714 610
rect 656 530 714 570
rect 656 490 668 530
rect 702 490 714 530
rect 656 450 714 490
rect 656 410 668 450
rect 702 410 714 450
rect 656 370 714 410
rect 656 330 668 370
rect 702 330 714 370
rect 656 290 714 330
rect 656 250 668 290
rect 702 250 714 290
rect 656 210 714 250
rect 656 172 668 210
rect 702 172 714 210
rect 656 156 714 172
rect 1074 982 1086 1015
rect 1492 1048 1550 1348
rect 2302 1298 2336 1338
rect 2302 1218 2336 1258
rect 2302 1138 2336 1178
rect 1120 982 1132 1015
rect 1074 942 1132 982
rect 1074 902 1086 942
rect 1120 902 1132 942
rect 1074 862 1132 902
rect 1074 822 1086 862
rect 1120 822 1132 862
rect 1074 782 1132 822
rect 1074 742 1086 782
rect 1120 742 1132 782
rect 1074 702 1132 742
rect 1074 662 1086 702
rect 1120 662 1132 702
rect 1074 622 1132 662
rect 1074 582 1086 622
rect 1120 582 1132 622
rect 1074 542 1132 582
rect 1074 502 1086 542
rect 1120 502 1132 542
rect 1074 462 1132 502
rect 1074 422 1086 462
rect 1120 422 1132 462
rect 1074 382 1132 422
rect 1074 342 1086 382
rect 1120 342 1132 382
rect 1074 302 1132 342
rect 1074 262 1086 302
rect 1120 262 1132 302
rect 1074 222 1132 262
rect 1074 172 1086 222
rect 1120 172 1132 222
rect 1074 96 1132 172
rect 1492 982 1504 1048
rect 1538 982 1550 1048
rect 1922 1048 1956 1064
rect 1492 942 1550 982
rect 1492 902 1504 942
rect 1538 902 1550 942
rect 1492 862 1550 902
rect 1492 822 1504 862
rect 1538 822 1550 862
rect 1492 782 1550 822
rect 1492 742 1504 782
rect 1538 742 1550 782
rect 1492 702 1550 742
rect 1492 662 1504 702
rect 1538 662 1550 702
rect 1492 622 1550 662
rect 1492 582 1504 622
rect 1538 582 1550 622
rect 1492 542 1550 582
rect 1492 502 1504 542
rect 1538 502 1550 542
rect 1492 462 1550 502
rect 1492 422 1504 462
rect 1538 422 1550 462
rect 1492 382 1550 422
rect 1492 342 1504 382
rect 1538 342 1550 382
rect 1492 302 1550 342
rect 1492 262 1504 302
rect 1538 262 1550 302
rect 1492 222 1550 262
rect 1492 172 1504 222
rect 1538 172 1550 222
rect 1492 156 1550 172
rect 1910 982 1922 1015
rect 2302 1058 2336 1098
rect 1956 1015 1961 1017
rect 1956 982 1968 1015
rect 1910 942 1968 982
rect 1910 902 1922 942
rect 1956 902 1968 942
rect 1910 862 1968 902
rect 1910 822 1922 862
rect 1956 822 1968 862
rect 1910 782 1968 822
rect 1910 742 1922 782
rect 1956 742 1968 782
rect 1910 702 1968 742
rect 1910 662 1922 702
rect 1956 662 1968 702
rect 1910 622 1968 662
rect 1910 582 1922 622
rect 1956 582 1968 622
rect 1910 542 1968 582
rect 2302 978 2336 1018
rect 2302 898 2336 938
rect 2302 818 2336 858
rect 2302 738 2336 778
rect 2302 658 2336 698
rect 2404 1552 2462 1606
rect 2404 1512 2416 1552
rect 2450 1512 2462 1552
rect 2404 1472 2462 1512
rect 2404 1432 2416 1472
rect 2450 1432 2462 1472
rect 2404 1392 2462 1432
rect 2404 1352 2416 1392
rect 2450 1352 2462 1392
rect 2404 1312 2462 1352
rect 2404 1272 2416 1312
rect 2450 1272 2462 1312
rect 2404 1232 2462 1272
rect 2404 1192 2416 1232
rect 2450 1192 2462 1232
rect 2404 1152 2462 1192
rect 2404 1112 2416 1152
rect 2450 1112 2462 1152
rect 2404 1072 2462 1112
rect 2404 1032 2416 1072
rect 2450 1032 2462 1072
rect 2404 992 2462 1032
rect 2404 952 2416 992
rect 2450 952 2462 992
rect 2404 912 2462 952
rect 2404 872 2416 912
rect 2450 872 2462 912
rect 2404 832 2462 872
rect 2404 792 2416 832
rect 2450 792 2462 832
rect 2404 752 2462 792
rect 2404 710 2416 752
rect 2450 710 2462 752
rect 2404 640 2462 710
rect 2822 1586 2880 1694
rect 2822 1544 2834 1586
rect 2868 1544 2880 1586
rect 2822 1504 2880 1544
rect 2822 1464 2834 1504
rect 2868 1464 2880 1504
rect 2822 1424 2880 1464
rect 2822 1384 2834 1424
rect 2868 1384 2880 1424
rect 2822 1344 2880 1384
rect 2822 1304 2834 1344
rect 2868 1304 2880 1344
rect 2822 1264 2880 1304
rect 2822 1224 2834 1264
rect 2868 1224 2880 1264
rect 2822 1184 2880 1224
rect 2822 1144 2834 1184
rect 2868 1144 2880 1184
rect 2822 1104 2880 1144
rect 2822 1064 2834 1104
rect 2868 1064 2880 1104
rect 2822 1024 2880 1064
rect 2822 984 2834 1024
rect 2868 984 2880 1024
rect 2822 944 2880 984
rect 2822 904 2834 944
rect 2868 904 2880 944
rect 2822 864 2880 904
rect 2822 824 2834 864
rect 2868 824 2880 864
rect 2822 784 2880 824
rect 2822 744 2834 784
rect 2868 744 2880 784
rect 2822 694 2880 744
rect 3240 1552 3298 1606
rect 3240 1512 3252 1552
rect 3286 1512 3298 1552
rect 3240 1472 3298 1512
rect 3240 1432 3252 1472
rect 3286 1432 3298 1472
rect 3240 1392 3298 1432
rect 3240 1352 3252 1392
rect 3286 1352 3298 1392
rect 3240 1312 3298 1352
rect 3240 1272 3252 1312
rect 3286 1272 3298 1312
rect 3240 1232 3298 1272
rect 3240 1192 3252 1232
rect 3286 1192 3298 1232
rect 3240 1152 3298 1192
rect 3240 1112 3252 1152
rect 3286 1112 3298 1152
rect 3240 1072 3298 1112
rect 3240 1032 3252 1072
rect 3286 1032 3298 1072
rect 3240 992 3298 1032
rect 3240 952 3252 992
rect 3286 952 3298 992
rect 3240 912 3298 952
rect 3240 872 3252 912
rect 3286 872 3298 912
rect 3240 832 3298 872
rect 3240 792 3252 832
rect 3286 792 3298 832
rect 3240 752 3298 792
rect 3240 710 3252 752
rect 3286 710 3298 752
rect 3240 640 3298 710
rect 3366 1532 3400 1560
rect 3880 1496 4120 1512
rect 3880 1472 3902 1496
rect 3366 1432 3400 1472
rect 3366 1352 3400 1392
rect 3780 1466 3902 1472
rect 3982 1466 4028 1496
rect 4108 1466 4120 1496
rect 3780 1348 3786 1466
rect 3876 1416 3902 1466
rect 3876 1382 3914 1416
rect 3876 1348 3902 1382
rect 3366 1272 3400 1312
rect 3880 1302 3902 1348
rect 3982 1302 4028 1348
rect 4108 1302 4120 1348
rect 3880 1286 4120 1302
rect 3366 1192 3400 1232
rect 3366 1112 3400 1152
rect 3366 1032 3400 1072
rect 3366 952 3400 992
rect 3366 872 3400 912
rect 3366 792 3400 832
rect 3366 712 3400 752
rect 3366 640 3400 659
rect 2336 634 2771 640
rect 2405 607 2443 634
rect 2527 607 2565 634
rect 2649 607 2687 634
rect 2931 634 3400 640
rect 3015 607 3053 634
rect 2405 573 2436 607
rect 2527 573 2536 607
rect 2656 573 2687 607
rect 2771 573 2776 607
rect 2816 573 2856 607
rect 2896 573 2931 607
rect 3015 573 3016 607
rect 2405 550 2443 573
rect 2527 550 2565 573
rect 2649 550 2687 573
rect 2302 544 2771 550
rect 3015 550 3053 573
rect 3137 550 3175 634
rect 3259 607 3297 634
rect 3259 550 3297 573
rect 2931 544 3400 550
rect 3833 950 3891 966
rect 3833 902 3845 950
rect 3879 902 3891 950
rect 3833 862 3891 902
rect 3833 822 3845 862
rect 3879 822 3891 862
rect 3833 782 3891 822
rect 3833 742 3845 782
rect 3879 742 3891 782
rect 3833 702 3891 742
rect 3833 662 3845 702
rect 3879 662 3891 702
rect 3833 622 3891 662
rect 3833 582 3845 622
rect 3879 582 3891 622
rect 1910 502 1922 542
rect 1956 502 1968 542
rect 1910 462 1968 502
rect 1910 422 1922 462
rect 1956 422 1968 462
rect 1910 382 1968 422
rect 1910 342 1922 382
rect 1956 342 1968 382
rect 1910 302 1968 342
rect 1910 262 1922 302
rect 1956 262 1968 302
rect 1910 222 1968 262
rect 1910 172 1922 222
rect 1956 172 1968 222
rect 1910 96 1968 172
rect 3833 542 3891 582
rect 3833 502 3845 542
rect 3879 502 3891 542
rect 3833 462 3891 502
rect 3833 422 3845 462
rect 3879 422 3891 462
rect 3833 382 3891 422
rect 3833 342 3845 382
rect 3879 342 3891 382
rect 3833 302 3891 342
rect 3833 262 3845 302
rect 3879 262 3891 302
rect 3833 222 3891 262
rect 3833 174 3845 222
rect 3879 174 3891 222
rect 3833 96 3891 174
rect 4250 950 4309 1694
rect 5127 1506 5186 2411
rect 5546 3187 5604 3264
rect 5546 3139 5558 3187
rect 5592 3139 5604 3187
rect 5546 3099 5604 3139
rect 5546 3059 5558 3099
rect 5592 3059 5604 3099
rect 5546 3019 5604 3059
rect 5546 2979 5558 3019
rect 5592 2979 5604 3019
rect 5546 2939 5604 2979
rect 5546 2899 5558 2939
rect 5592 2899 5604 2939
rect 5546 2859 5604 2899
rect 5546 2819 5558 2859
rect 5592 2819 5604 2859
rect 5546 2779 5604 2819
rect 5546 2739 5558 2779
rect 5592 2739 5604 2779
rect 5546 2699 5604 2739
rect 5546 2659 5558 2699
rect 5592 2659 5604 2699
rect 5546 2619 5604 2659
rect 5546 2579 5558 2619
rect 5592 2579 5604 2619
rect 5546 2539 5604 2579
rect 5546 2499 5558 2539
rect 5592 2499 5604 2539
rect 5546 2459 5604 2499
rect 5546 2411 5558 2459
rect 5592 2411 5604 2459
rect 5546 2395 5604 2411
rect 5310 2060 5546 2068
rect 5310 1858 5326 2060
rect 5406 2002 5446 2060
rect 5526 2012 5546 2060
rect 5526 2002 5646 2012
rect 5526 1972 5556 2002
rect 5516 1938 5556 1972
rect 5526 1902 5556 1938
rect 5636 1902 5646 2002
rect 5406 1858 5446 1902
rect 5526 1892 5646 1902
rect 5526 1858 5546 1892
rect 5310 1852 5546 1858
rect 5127 1485 5140 1506
rect 5081 1479 5140 1485
rect 5174 1485 5186 1506
rect 5546 1506 5604 1522
rect 5174 1479 5229 1485
rect 5081 1335 5093 1479
rect 5217 1335 5229 1479
rect 5081 1329 5140 1335
rect 5127 1302 5140 1329
rect 5174 1329 5229 1335
rect 5546 1462 5558 1506
rect 5592 1462 5604 1506
rect 5546 1422 5604 1462
rect 5546 1382 5558 1422
rect 5592 1382 5604 1422
rect 5546 1342 5604 1382
rect 5174 1302 5186 1329
rect 5127 1262 5186 1302
rect 5127 1222 5140 1262
rect 5174 1222 5186 1262
rect 5026 1172 5060 1212
rect 5026 1092 5060 1132
rect 5026 1012 5060 1052
rect 4250 902 4263 950
rect 4297 902 4309 950
rect 4250 862 4309 902
rect 4250 822 4263 862
rect 4297 822 4309 862
rect 4250 782 4309 822
rect 4250 742 4263 782
rect 4297 742 4309 782
rect 4250 702 4309 742
rect 4250 662 4263 702
rect 4297 662 4309 702
rect 4250 622 4309 662
rect 4250 582 4263 622
rect 4297 582 4309 622
rect 4250 542 4309 582
rect 4250 502 4263 542
rect 4297 502 4309 542
rect 4250 462 4309 502
rect 4250 422 4263 462
rect 4297 422 4309 462
rect 4250 382 4309 422
rect 4250 342 4263 382
rect 4297 342 4309 382
rect 4250 302 4309 342
rect 4250 262 4263 302
rect 4297 262 4309 302
rect 4250 222 4309 262
rect 4250 174 4263 222
rect 4297 174 4309 222
rect 4250 158 4309 174
rect 4669 950 4727 966
rect 4669 902 4681 950
rect 4715 902 4727 950
rect 4669 862 4727 902
rect 4669 822 4681 862
rect 4715 822 4727 862
rect 4669 782 4727 822
rect 4669 742 4681 782
rect 4715 742 4727 782
rect 4669 702 4727 742
rect 4669 662 4681 702
rect 4715 662 4727 702
rect 4669 622 4727 662
rect 4669 582 4681 622
rect 4715 582 4727 622
rect 5026 932 5060 972
rect 5026 852 5060 892
rect 5026 772 5060 812
rect 5026 692 5060 732
rect 5127 1182 5186 1222
rect 5127 1142 5140 1182
rect 5174 1142 5186 1182
rect 5127 1102 5186 1142
rect 5127 1062 5140 1102
rect 5174 1062 5186 1102
rect 5127 1022 5186 1062
rect 5127 982 5140 1022
rect 5174 982 5186 1022
rect 5127 942 5186 982
rect 5127 902 5140 942
rect 5174 902 5186 942
rect 5127 862 5186 902
rect 5127 822 5140 862
rect 5174 822 5186 862
rect 5127 782 5186 822
rect 5127 730 5140 782
rect 5174 730 5186 782
rect 5127 714 5186 730
rect 5546 1302 5558 1342
rect 5592 1302 5604 1342
rect 5546 1262 5604 1302
rect 5546 1222 5558 1262
rect 5592 1222 5604 1262
rect 5546 1182 5604 1222
rect 5546 1142 5558 1182
rect 5592 1142 5604 1182
rect 5546 1102 5604 1142
rect 5546 1062 5558 1102
rect 5592 1062 5604 1102
rect 5546 1022 5604 1062
rect 5546 982 5558 1022
rect 5592 982 5604 1022
rect 5546 942 5604 982
rect 5546 902 5558 942
rect 5592 902 5604 942
rect 5546 862 5604 902
rect 5546 822 5558 862
rect 5592 822 5604 862
rect 5546 782 5604 822
rect 5546 730 5558 782
rect 5592 730 5604 782
rect 5026 583 5060 652
rect 5546 640 5604 730
rect 5672 1493 5706 1523
rect 5672 1410 5706 1450
rect 5672 1330 5706 1370
rect 5672 1250 5706 1290
rect 5672 1170 5706 1210
rect 5672 1090 5706 1130
rect 5672 1010 5706 1050
rect 5672 930 5706 970
rect 5672 850 5706 890
rect 5672 770 5706 810
rect 5672 690 5706 730
rect 5287 634 5672 640
rect 5340 617 5378 634
rect 5462 617 5500 634
rect 5584 617 5622 634
rect 5120 583 5160 617
rect 5200 583 5240 617
rect 5360 583 5378 617
rect 5462 583 5480 617
rect 5610 583 5622 617
rect 4669 542 4727 582
rect 5340 550 5378 583
rect 5462 550 5500 583
rect 5584 550 5622 583
rect 5287 544 5706 550
rect 4669 502 4681 542
rect 4715 502 4727 542
rect 4669 462 4727 502
rect 4669 422 4681 462
rect 4715 422 4727 462
rect 4669 382 4727 422
rect 4669 342 4681 382
rect 4715 342 4727 382
rect 4669 302 4727 342
rect 4669 262 4681 302
rect 4715 262 4727 302
rect 4669 222 4727 262
rect 4669 174 4681 222
rect 4715 174 4727 222
rect 4669 96 4727 174
rect 136 90 605 96
rect 239 6 277 90
rect 361 6 399 90
rect 483 6 521 90
rect 136 0 605 6
rect 818 90 1390 96
rect 902 6 940 90
rect 1024 6 1062 90
rect 1146 6 1184 90
rect 1268 6 1306 90
rect 818 0 1390 6
rect 1601 90 2070 96
rect 1685 6 1723 90
rect 1807 6 1845 90
rect 1929 6 1967 90
rect 1601 0 2070 6
rect 3731 90 4200 96
rect 3815 6 3853 90
rect 3937 6 3975 90
rect 4059 6 4097 90
rect 3731 0 4200 6
rect 4360 90 4829 96
rect 4463 6 4501 90
rect 4585 6 4623 90
rect 4707 6 4745 90
rect 4360 0 4829 6
<< viali >>
rect 1466 3270 1569 3354
rect 1607 3270 1691 3354
rect 1729 3270 1813 3354
rect 1851 3270 1935 3354
rect 2146 3270 2230 3354
rect 2268 3270 2352 3354
rect 2390 3270 2474 3354
rect 2512 3270 2596 3354
rect 2634 3270 2718 3354
rect 2931 3270 3015 3354
rect 3053 3270 3137 3354
rect 3175 3270 3259 3354
rect 3297 3270 3400 3354
rect 4608 3270 4710 3354
rect 4750 3270 4832 3354
rect 4872 3270 4954 3354
rect 4994 3270 5077 3354
rect 5237 3270 5321 3354
rect 5359 3270 5443 3354
rect 5481 3270 5565 3354
rect 5603 3270 5706 3354
rect 136 2779 239 2810
rect 277 2779 361 2810
rect 136 2745 232 2779
rect 232 2745 239 2779
rect 277 2745 280 2779
rect 280 2745 320 2779
rect 320 2745 360 2779
rect 360 2745 361 2779
rect 136 2726 239 2745
rect 277 2726 361 2745
rect 399 2779 483 2810
rect 521 2779 605 2810
rect 801 2779 885 2810
rect 923 2779 1007 2810
rect 1045 2779 1129 2810
rect 399 2745 400 2779
rect 400 2745 440 2779
rect 440 2745 480 2779
rect 480 2745 483 2779
rect 521 2745 560 2779
rect 560 2745 600 2779
rect 600 2745 605 2779
rect 801 2745 840 2779
rect 840 2745 880 2779
rect 880 2745 885 2779
rect 923 2745 960 2779
rect 960 2745 1000 2779
rect 1000 2745 1007 2779
rect 1045 2745 1100 2779
rect 1100 2745 1129 2779
rect 399 2726 483 2745
rect 521 2726 605 2745
rect 801 2726 885 2745
rect 923 2726 1007 2745
rect 1045 2726 1129 2745
rect 1167 2726 1270 2810
rect 286 1426 296 1500
rect 296 1426 376 1500
rect 376 1426 410 1500
rect 410 1426 488 1500
rect 286 1390 488 1426
rect 286 1312 296 1390
rect 296 1312 376 1390
rect 376 1312 410 1390
rect 410 1312 488 1390
rect 3731 2730 3815 2810
rect 3853 2778 3937 2810
rect 3975 2778 4059 2810
rect 4097 2778 4181 2810
rect 3853 2744 3880 2778
rect 3880 2744 3920 2778
rect 3920 2744 3937 2778
rect 3975 2744 4000 2778
rect 4000 2744 4040 2778
rect 4040 2744 4059 2778
rect 4097 2744 4120 2778
rect 4120 2744 4160 2778
rect 4160 2744 4181 2778
rect 3731 2726 3765 2730
rect 3765 2726 3815 2730
rect 3853 2726 3937 2744
rect 3975 2726 4059 2744
rect 4097 2726 4181 2744
rect 3080 2000 3220 2018
rect 2600 1880 2616 2000
rect 2616 1880 2720 2000
rect 2760 1880 2776 2000
rect 2776 1880 2880 2000
rect 2920 1880 2936 2000
rect 2936 1880 3040 2000
rect 3080 1880 3096 2000
rect 3096 1880 3216 2000
rect 3216 1880 3220 2000
rect 3260 1892 3388 2018
rect 4713 1892 4813 2012
rect 1492 1348 1656 1468
rect 3786 1348 3876 1466
rect 3914 1416 3982 1466
rect 3982 1416 4028 1466
rect 4028 1416 4108 1466
rect 4108 1416 4120 1466
rect 3914 1382 4120 1416
rect 3914 1348 3982 1382
rect 3982 1348 4028 1382
rect 4028 1348 4108 1382
rect 4108 1348 4120 1382
rect 2302 624 2336 634
rect 2336 624 2405 634
rect 2302 550 2405 624
rect 2443 607 2527 634
rect 2565 607 2649 634
rect 2687 607 2771 634
rect 2931 607 3015 634
rect 3053 607 3137 634
rect 2443 573 2496 607
rect 2496 573 2527 607
rect 2565 573 2576 607
rect 2576 573 2616 607
rect 2616 573 2649 607
rect 2687 573 2696 607
rect 2696 573 2736 607
rect 2736 573 2771 607
rect 2931 573 2936 607
rect 2936 573 2976 607
rect 2976 573 3015 607
rect 3053 573 3056 607
rect 3056 573 3096 607
rect 3096 573 3136 607
rect 3136 573 3137 607
rect 2443 550 2527 573
rect 2565 550 2649 573
rect 2687 550 2771 573
rect 2931 550 3015 573
rect 3053 550 3137 573
rect 3175 607 3259 634
rect 3297 607 3400 634
rect 3175 573 3176 607
rect 3176 573 3216 607
rect 3216 573 3256 607
rect 3256 573 3259 607
rect 3297 573 3304 607
rect 3304 573 3400 607
rect 3175 550 3259 573
rect 3297 550 3400 573
rect 5326 1972 5406 2002
rect 5406 1972 5446 2002
rect 5446 1972 5516 2002
rect 5326 1938 5516 1972
rect 5326 1902 5406 1938
rect 5406 1902 5446 1938
rect 5446 1902 5516 1938
rect 5556 1902 5636 2002
rect 5093 1462 5140 1479
rect 5140 1462 5174 1479
rect 5174 1462 5217 1479
rect 5093 1422 5217 1462
rect 5093 1382 5140 1422
rect 5140 1382 5174 1422
rect 5174 1382 5217 1422
rect 5093 1342 5217 1382
rect 5093 1335 5140 1342
rect 5140 1335 5174 1342
rect 5174 1335 5217 1342
rect 5256 617 5340 634
rect 5378 617 5462 634
rect 5500 617 5584 634
rect 5622 631 5672 634
rect 5672 631 5706 634
rect 5256 583 5280 617
rect 5280 583 5320 617
rect 5320 583 5340 617
rect 5378 583 5400 617
rect 5400 583 5440 617
rect 5440 583 5462 617
rect 5500 583 5520 617
rect 5520 583 5560 617
rect 5560 583 5584 617
rect 5256 550 5340 583
rect 5378 550 5462 583
rect 5500 550 5584 583
rect 5622 550 5706 631
rect 136 6 239 90
rect 277 6 361 90
rect 399 6 483 90
rect 521 6 605 90
rect 818 6 902 90
rect 940 6 1024 90
rect 1062 6 1146 90
rect 1184 6 1268 90
rect 1306 6 1390 90
rect 1601 6 1685 90
rect 1723 6 1807 90
rect 1845 6 1929 90
rect 1967 6 2070 90
rect 3731 6 3815 90
rect 3853 6 3937 90
rect 3975 6 4059 90
rect 4097 6 4200 90
rect 4360 6 4463 90
rect 4501 6 4585 90
rect 4623 6 4707 90
rect 4745 6 4829 90
<< metal1 >>
rect 0 3354 5900 3360
rect 0 3270 1466 3354
rect 1569 3270 1607 3354
rect 1691 3270 1729 3354
rect 1813 3270 1851 3354
rect 1935 3270 2146 3354
rect 2230 3270 2268 3354
rect 2352 3270 2390 3354
rect 2474 3270 2512 3354
rect 2596 3270 2634 3354
rect 2718 3270 2931 3354
rect 3015 3270 3053 3354
rect 3137 3270 3175 3354
rect 3259 3270 3297 3354
rect 3400 3270 4608 3354
rect 4710 3270 4750 3354
rect 4832 3270 4872 3354
rect 4954 3270 4994 3354
rect 5077 3270 5237 3354
rect 5321 3270 5359 3354
rect 5443 3270 5481 3354
rect 5565 3270 5603 3354
rect 5706 3270 5900 3354
rect 0 3264 5900 3270
rect 0 2810 5900 2816
rect 0 2726 136 2810
rect 239 2726 277 2810
rect 361 2726 399 2810
rect 483 2726 521 2810
rect 605 2726 801 2810
rect 885 2726 923 2810
rect 1007 2726 1045 2810
rect 1129 2726 1167 2810
rect 1270 2726 3731 2810
rect 3815 2726 3853 2810
rect 3937 2726 3975 2810
rect 4059 2726 4097 2810
rect 4181 2726 5900 2810
rect 0 2720 5900 2726
rect 2580 2018 3400 2024
rect 2580 2012 3080 2018
rect 0 2000 3080 2012
rect 0 1892 2600 2000
rect 2580 1880 2600 1892
rect 2720 1880 2760 2000
rect 2880 1880 2920 2000
rect 3040 1880 3080 2000
rect 3220 1892 3260 2018
rect 3388 1892 3400 2018
rect 3220 1880 3400 1892
rect 4707 2012 4819 2024
rect 4707 1892 4713 2012
rect 4813 2002 5900 2012
rect 4813 1902 5326 2002
rect 5516 1902 5556 2002
rect 5636 1902 5900 2002
rect 4813 1892 5900 1902
rect 4707 1880 4819 1892
rect 2580 1874 3240 1880
rect 280 1500 506 1516
rect 280 1473 286 1500
rect 0 1341 286 1473
rect 280 1312 286 1341
rect 488 1312 506 1500
rect 5081 1479 5229 1485
rect 1480 1473 4132 1474
rect 5081 1473 5093 1479
rect 1480 1468 5093 1473
rect 1480 1348 1492 1468
rect 1656 1466 5093 1468
rect 1656 1348 3786 1466
rect 3876 1348 3914 1466
rect 4120 1348 5093 1466
rect 1480 1342 5093 1348
rect 3434 1341 5093 1342
rect 5081 1335 5093 1341
rect 5217 1473 5229 1479
rect 5217 1341 5900 1473
rect 5217 1335 5229 1341
rect 5081 1329 5229 1335
rect 280 1296 506 1312
rect 0 634 5900 640
rect 0 550 2302 634
rect 2405 550 2443 634
rect 2527 550 2565 634
rect 2649 550 2687 634
rect 2771 550 2931 634
rect 3015 550 3053 634
rect 3137 550 3175 634
rect 3259 550 3297 634
rect 3400 550 5256 634
rect 5340 550 5378 634
rect 5462 550 5500 634
rect 5584 550 5622 634
rect 5706 550 5900 634
rect 0 544 5900 550
rect 0 90 5900 96
rect 0 6 136 90
rect 239 6 277 90
rect 361 6 399 90
rect 483 6 521 90
rect 605 6 818 90
rect 902 6 940 90
rect 1024 6 1062 90
rect 1146 6 1184 90
rect 1268 6 1306 90
rect 1390 6 1601 90
rect 1685 6 1723 90
rect 1807 6 1845 90
rect 1929 6 1967 90
rect 2070 6 3731 90
rect 3815 6 3853 90
rect 3937 6 3975 90
rect 4059 6 4097 90
rect 4200 6 4360 90
rect 4463 6 4501 90
rect 4585 6 4623 90
rect 4707 6 4745 90
rect 4829 6 5900 90
rect 0 0 5900 6
<< labels >>
flabel metal1 2376 2720 2776 2804 1 FreeSans 400 0 0 0 vdd
flabel metal1 2336 3276 2736 3360 1 FreeSans 400 0 0 0 vss
flabel metal1 800 558 1200 642 5 FreeSans 400 180 0 0 vdd
flabel metal1 2292 0 2844 96 1 FreeSans 400 0 0 0 vss
flabel metal1 5241 1346 5341 1466 1 FreeSans 400 1 0 0 outn
flabel metal1 4819 1892 4919 2012 1 FreeSans 400 1 0 0 outp
flabel metal1 174 1347 274 1467 1 FreeSans 400 1 0 0 inn
flabel metal1 1600 1892 1700 2012 1 FreeSans 400 1 0 0 inp
<< end >>
