magic
tech sky130A
timestamp 1637571367
<< nwell >>
rect 0 0 225 450
<< pdiff >>
rect 47 387 153 404
rect 47 369 51 387
rect 69 369 91 387
rect 109 369 131 387
rect 149 369 153 387
rect 47 359 153 369
rect 48 356 152 359
rect 49 353 151 356
rect 50 350 150 353
rect 50 97 150 100
rect 49 94 151 97
rect 48 91 152 94
rect 47 81 153 91
rect 47 63 51 81
rect 69 63 91 81
rect 109 63 131 81
rect 149 63 153 81
rect 47 46 153 63
<< pdiffc >>
rect 51 369 69 387
rect 91 369 109 387
rect 131 369 149 387
rect 51 63 69 81
rect 91 63 109 81
rect 131 63 149 81
<< nsubdiff >>
rect 180 232 200 244
rect 180 200 200 212
<< nsubdiffcont >>
rect 180 212 200 232
<< pdiffres >>
rect 50 100 150 350
<< locali >>
rect 46 388 154 397
rect 46 368 50 388
rect 70 368 90 388
rect 110 368 130 388
rect 150 368 154 388
rect 46 359 154 368
rect 180 232 200 241
rect 180 203 200 212
rect 46 82 154 91
rect 46 62 50 82
rect 70 62 90 82
rect 110 62 130 82
rect 150 62 154 82
rect 46 53 154 62
<< viali >>
rect 50 387 70 388
rect 50 369 51 387
rect 51 369 69 387
rect 69 369 70 387
rect 50 368 70 369
rect 90 387 110 388
rect 90 369 91 387
rect 91 369 109 387
rect 109 369 110 387
rect 90 368 110 369
rect 130 387 150 388
rect 130 369 131 387
rect 131 369 149 387
rect 149 369 150 387
rect 130 368 150 369
rect 50 81 70 82
rect 50 63 51 81
rect 51 63 69 81
rect 69 63 70 81
rect 50 62 70 63
rect 90 81 110 82
rect 90 63 91 81
rect 91 63 109 81
rect 109 63 110 81
rect 90 62 110 63
rect 130 81 150 82
rect 130 63 131 81
rect 131 63 149 81
rect 149 63 150 81
rect 130 62 150 63
<< metal1 >>
rect 46 388 154 397
rect 46 368 50 388
rect 70 368 90 388
rect 110 368 130 388
rect 150 368 154 388
rect 46 359 154 368
rect 46 85 154 91
rect 46 59 47 85
rect 73 59 87 85
rect 113 59 127 85
rect 153 59 154 85
rect 46 53 154 59
<< via1 >>
rect 47 82 73 85
rect 47 62 50 82
rect 50 62 70 82
rect 70 62 73 82
rect 47 59 73 62
rect 87 82 113 85
rect 87 62 90 82
rect 90 62 110 82
rect 110 62 113 82
rect 87 59 113 62
rect 127 82 153 85
rect 127 62 130 82
rect 130 62 150 82
rect 150 62 153 82
rect 127 59 153 62
<< metal2 >>
rect 41 86 159 91
rect 41 58 46 86
rect 74 58 86 86
rect 114 58 126 86
rect 154 58 159 86
rect 41 53 159 58
<< via2 >>
rect 46 85 74 86
rect 46 59 47 85
rect 47 59 73 85
rect 73 59 74 85
rect 46 58 74 59
rect 86 85 114 86
rect 86 59 87 85
rect 87 59 113 85
rect 113 59 114 85
rect 86 58 114 59
rect 126 85 154 86
rect 126 59 127 85
rect 127 59 153 85
rect 153 59 154 85
rect 126 58 154 59
<< metal3 >>
rect 41 86 159 91
rect 41 58 46 86
rect 74 58 86 86
rect 114 58 126 86
rect 154 58 159 86
rect 41 53 159 58
<< end >>
