magic
tech sky130A
magscale 1 2
timestamp 1637949574
<< nwell >>
rect -200 5142 336 5190
rect 599 5142 951 5190
rect -162 5120 38 5142
rect 599 5120 865 5142
<< nsubdiff >>
rect -162 5120 -119 5154
rect -85 5120 -39 5154
rect -5 5120 38 5154
rect 637 5120 680 5154
rect 714 5120 760 5154
rect 794 5120 837 5154
<< nsubdiffcont >>
rect -119 5120 -85 5154
rect -39 5120 -5 5154
rect 680 5120 714 5154
rect 760 5120 794 5154
<< poly >>
rect 20500 3900 20600 3973
rect 20500 3872 20673 3900
rect 20500 3838 20538 3872
rect 20572 3838 20673 3872
rect 20500 3800 20673 3838
<< polycont >>
rect 20538 3838 20572 3872
<< locali >>
rect -162 5120 -119 5154
rect -85 5120 -39 5154
rect -5 5120 38 5154
rect 637 5120 680 5154
rect 714 5120 760 5154
rect 794 5121 837 5154
rect 794 5120 850 5121
rect 336 4950 601 4992
rect 281 4948 601 4950
rect 281 4906 380 4948
rect 557 4907 601 4948
rect 557 4863 654 4907
rect 442 4849 502 4862
rect 442 4815 455 4849
rect 489 4815 502 4849
rect 442 4696 502 4815
rect 20220 4857 20280 4870
rect 20220 4823 20233 4857
rect 20267 4823 20280 4857
rect 20220 4810 20280 4823
rect 20320 4857 20380 4870
rect 20320 4823 20333 4857
rect 20367 4823 20380 4857
rect 20320 4810 20380 4823
rect 20420 4857 20480 4870
rect 20420 4823 20433 4857
rect 20467 4823 20480 4857
rect 20420 4810 20480 4823
rect 20520 4857 20580 4870
rect 20520 4823 20533 4857
rect 20567 4823 20580 4857
rect 20520 4810 20580 4823
rect 281 4636 502 4696
rect 20400 3900 20600 3973
rect 20400 3872 20673 3900
rect 20400 3871 20538 3872
rect 20400 3837 20431 3871
rect 20465 3837 20535 3871
rect 20572 3838 20673 3872
rect 20569 3837 20673 3838
rect 20400 3767 20673 3837
rect 20400 3733 20431 3767
rect 20465 3733 20535 3767
rect 20569 3733 20673 3767
rect 20400 3700 20673 3733
rect 21504 3875 21700 3900
rect 21504 3820 21519 3875
rect 21521 3867 21700 3875
rect 21521 3833 21534 3867
rect 21568 3833 21632 3867
rect 21666 3833 21700 3867
rect 21521 3820 21700 3833
rect 21504 3767 21700 3820
rect 21504 3733 21534 3767
rect 21568 3733 21632 3767
rect 21666 3733 21700 3767
rect 21504 3700 21700 3733
<< viali >>
rect 455 4815 489 4849
rect 20233 4823 20267 4857
rect 20333 4823 20367 4857
rect 20433 4823 20467 4857
rect 20533 4823 20567 4857
rect 20431 3837 20465 3871
rect 20535 3838 20538 3871
rect 20538 3838 20569 3871
rect 20535 3837 20569 3838
rect 20431 3733 20465 3767
rect 20535 3733 20569 3767
rect 21534 3833 21568 3867
rect 21632 3833 21666 3867
rect 21534 3733 21568 3767
rect 21632 3733 21666 3767
<< metal1 >>
rect 1680 5854 1914 5950
rect -200 5120 865 5152
rect -200 5056 640 5120
rect 436 4849 1698 4862
rect 436 4815 455 4849
rect 489 4815 1698 4849
rect 436 4802 1698 4815
rect 1152 4790 1698 4802
rect 5254 4790 5326 4862
rect 12334 4790 12406 4862
rect 15878 4790 15950 4862
rect 19508 4790 19622 4862
rect 19810 4790 20044 4862
rect 20200 4857 20601 4876
rect 20200 4823 20233 4857
rect 20267 4823 20333 4857
rect 20367 4823 20433 4857
rect 20467 4823 20533 4857
rect 20567 4823 20601 4857
rect 20200 4803 20601 4823
rect -200 4512 637 4608
rect 1152 3472 1224 4790
rect -502 3400 1224 3472
rect 1424 4246 1702 4318
rect 5254 4246 5326 4318
rect 8798 4246 8870 4318
rect 12334 4246 12406 4318
rect 15878 4246 15950 4318
rect 19504 4246 19772 4318
rect -502 1178 -430 3400
rect 1424 3200 1496 4246
rect -230 3128 1496 3200
rect 2400 3206 2600 3230
rect 2452 3154 2474 3206
rect 2526 3154 2548 3206
rect 2400 3134 2600 3154
rect 3600 3206 3800 3230
rect 3652 3154 3674 3206
rect 3726 3154 3748 3206
rect 3600 3134 3800 3154
rect 4800 3206 5000 3230
rect 4852 3154 4874 3206
rect 4926 3154 4948 3206
rect 4800 3134 5000 3154
rect 6000 3206 6200 3230
rect 6052 3154 6074 3206
rect 6126 3154 6148 3206
rect 6000 3134 6200 3154
rect 7200 3206 7400 3230
rect 7252 3154 7274 3206
rect 7326 3154 7348 3206
rect 7200 3134 7400 3154
rect 8400 3206 8600 3230
rect 8452 3154 8474 3206
rect 8526 3154 8548 3206
rect 8400 3134 8600 3154
rect 9600 3206 9800 3230
rect 9652 3154 9674 3206
rect 9726 3154 9748 3206
rect 9600 3134 9800 3154
rect 10800 3206 11000 3230
rect 10852 3154 10874 3206
rect 10926 3154 10948 3206
rect 10800 3134 11000 3154
rect 12000 3206 12200 3230
rect 12052 3154 12074 3206
rect 12126 3154 12148 3206
rect 12000 3134 12200 3154
rect 13200 3206 13400 3230
rect 13252 3154 13274 3206
rect 13326 3154 13348 3206
rect 13200 3134 13400 3154
rect 14400 3206 14600 3230
rect 14452 3154 14474 3206
rect 14526 3154 14548 3206
rect 14400 3134 14600 3154
rect 15600 3206 15800 3230
rect 15652 3154 15674 3206
rect 15726 3154 15748 3206
rect 15600 3134 15800 3154
rect 16800 3206 17000 3230
rect 16852 3154 16874 3206
rect 16926 3154 16948 3206
rect 16800 3134 17000 3154
rect 18000 3206 18200 3230
rect 18052 3154 18074 3206
rect 18126 3154 18148 3206
rect 18000 3134 18200 3154
rect 19200 3206 19400 3230
rect 19252 3154 19274 3206
rect 19326 3154 19348 3206
rect 19200 3134 19400 3154
rect 19700 3200 19772 4246
rect 19972 3472 20044 4790
rect 20400 3880 20600 3903
rect 20400 3828 20422 3880
rect 20474 3828 20526 3880
rect 20578 3828 20600 3880
rect 20400 3776 20600 3828
rect 20400 3724 20422 3776
rect 20474 3724 20526 3776
rect 20578 3724 20600 3776
rect 20400 3700 20600 3724
rect 21503 3876 21700 3900
rect 21503 3824 21525 3876
rect 21577 3824 21623 3876
rect 21675 3824 21700 3876
rect 21503 3776 21700 3824
rect 21503 3724 21525 3776
rect 21577 3724 21623 3776
rect 21675 3724 21700 3776
rect 21503 3700 21700 3724
rect 19972 3400 21872 3472
rect 19700 3128 21600 3200
rect -230 1722 -158 3128
rect 0 2810 200 2834
rect 52 2758 74 2810
rect 126 2758 148 2810
rect 0 2738 200 2758
rect 1200 2810 1400 2834
rect 1252 2758 1274 2810
rect 1326 2758 1348 2810
rect 1200 2738 1400 2758
rect 2400 2810 2600 2834
rect 2452 2758 2474 2810
rect 2526 2758 2548 2810
rect 2400 2738 2600 2758
rect 3600 2810 3800 2834
rect 3652 2758 3674 2810
rect 3726 2758 3748 2810
rect 3600 2738 3800 2758
rect 4800 2810 5000 2834
rect 4852 2758 4874 2810
rect 4926 2758 4948 2810
rect 4800 2738 5000 2758
rect 6000 2810 6200 2834
rect 6052 2758 6074 2810
rect 6126 2758 6148 2810
rect 6000 2738 6200 2758
rect 7200 2810 7400 2834
rect 7252 2758 7274 2810
rect 7326 2758 7348 2810
rect 7200 2738 7400 2758
rect 8400 2810 8600 2834
rect 8452 2758 8474 2810
rect 8526 2758 8548 2810
rect 8400 2738 8600 2758
rect 9600 2810 9800 2834
rect 9652 2758 9674 2810
rect 9726 2758 9748 2810
rect 9600 2738 9800 2758
rect 10800 2810 11000 2834
rect 10852 2758 10874 2810
rect 10926 2758 10948 2810
rect 10800 2738 11000 2758
rect 12000 2810 12200 2834
rect 12052 2758 12074 2810
rect 12126 2758 12148 2810
rect 12000 2738 12200 2758
rect 13200 2810 13400 2834
rect 13252 2758 13274 2810
rect 13326 2758 13348 2810
rect 13200 2738 13400 2758
rect 14400 2810 14600 2834
rect 14452 2758 14474 2810
rect 14526 2758 14548 2810
rect 14400 2738 14600 2758
rect 15600 2810 15800 2834
rect 15652 2758 15674 2810
rect 15726 2758 15748 2810
rect 15600 2738 15800 2758
rect 16800 2810 17000 2834
rect 16852 2758 16874 2810
rect 16926 2758 16948 2810
rect 16800 2738 17000 2758
rect 18000 2810 18200 2834
rect 18052 2758 18074 2810
rect 18126 2758 18148 2810
rect 18000 2738 18200 2758
rect 19200 2810 19400 2834
rect 19252 2758 19274 2810
rect 19326 2758 19348 2810
rect 19200 2738 19400 2758
rect 20400 2810 20600 2834
rect 20452 2758 20474 2810
rect 20526 2758 20548 2810
rect 20400 2738 20600 2758
rect 21156 2810 21356 2834
rect 21208 2758 21230 2810
rect 21282 2758 21304 2810
rect 21156 2738 21356 2758
rect 21528 1722 21600 3128
rect -230 1650 0 1722
rect 3554 1650 3626 1722
rect 7104 1650 7176 1722
rect 10634 1650 10706 1722
rect 14182 1650 14254 1722
rect 17728 1650 17800 1722
rect 21267 1650 21600 1722
rect 21800 1178 21872 3400
rect -502 1106 -130 1178
rect 10650 1106 10722 1178
rect 14182 1106 14254 1178
rect 21356 1106 21872 1178
<< via1 >>
rect 2400 3154 2452 3206
rect 2474 3154 2526 3206
rect 2548 3154 2600 3206
rect 3600 3154 3652 3206
rect 3674 3154 3726 3206
rect 3748 3154 3800 3206
rect 4800 3154 4852 3206
rect 4874 3154 4926 3206
rect 4948 3154 5000 3206
rect 6000 3154 6052 3206
rect 6074 3154 6126 3206
rect 6148 3154 6200 3206
rect 7200 3154 7252 3206
rect 7274 3154 7326 3206
rect 7348 3154 7400 3206
rect 8400 3154 8452 3206
rect 8474 3154 8526 3206
rect 8548 3154 8600 3206
rect 9600 3154 9652 3206
rect 9674 3154 9726 3206
rect 9748 3154 9800 3206
rect 10800 3154 10852 3206
rect 10874 3154 10926 3206
rect 10948 3154 11000 3206
rect 12000 3154 12052 3206
rect 12074 3154 12126 3206
rect 12148 3154 12200 3206
rect 13200 3154 13252 3206
rect 13274 3154 13326 3206
rect 13348 3154 13400 3206
rect 14400 3154 14452 3206
rect 14474 3154 14526 3206
rect 14548 3154 14600 3206
rect 15600 3154 15652 3206
rect 15674 3154 15726 3206
rect 15748 3154 15800 3206
rect 16800 3154 16852 3206
rect 16874 3154 16926 3206
rect 16948 3154 17000 3206
rect 18000 3154 18052 3206
rect 18074 3154 18126 3206
rect 18148 3154 18200 3206
rect 19200 3154 19252 3206
rect 19274 3154 19326 3206
rect 19348 3154 19400 3206
rect 20422 3871 20474 3880
rect 20422 3837 20431 3871
rect 20431 3837 20465 3871
rect 20465 3837 20474 3871
rect 20422 3828 20474 3837
rect 20526 3871 20578 3880
rect 20526 3837 20535 3871
rect 20535 3837 20569 3871
rect 20569 3837 20578 3871
rect 20526 3828 20578 3837
rect 20422 3767 20474 3776
rect 20422 3733 20431 3767
rect 20431 3733 20465 3767
rect 20465 3733 20474 3767
rect 20422 3724 20474 3733
rect 20526 3767 20578 3776
rect 20526 3733 20535 3767
rect 20535 3733 20569 3767
rect 20569 3733 20578 3767
rect 20526 3724 20578 3733
rect 21525 3867 21577 3876
rect 21525 3833 21534 3867
rect 21534 3833 21568 3867
rect 21568 3833 21577 3867
rect 21525 3824 21577 3833
rect 21623 3867 21675 3876
rect 21623 3833 21632 3867
rect 21632 3833 21666 3867
rect 21666 3833 21675 3867
rect 21623 3824 21675 3833
rect 21525 3767 21577 3776
rect 21525 3733 21534 3767
rect 21534 3733 21568 3767
rect 21568 3733 21577 3767
rect 21525 3724 21577 3733
rect 21623 3767 21675 3776
rect 21623 3733 21632 3767
rect 21632 3733 21666 3767
rect 21666 3733 21675 3767
rect 21623 3724 21675 3733
rect 0 2758 52 2810
rect 74 2758 126 2810
rect 148 2758 200 2810
rect 1200 2758 1252 2810
rect 1274 2758 1326 2810
rect 1348 2758 1400 2810
rect 2400 2758 2452 2810
rect 2474 2758 2526 2810
rect 2548 2758 2600 2810
rect 3600 2758 3652 2810
rect 3674 2758 3726 2810
rect 3748 2758 3800 2810
rect 4800 2758 4852 2810
rect 4874 2758 4926 2810
rect 4948 2758 5000 2810
rect 6000 2758 6052 2810
rect 6074 2758 6126 2810
rect 6148 2758 6200 2810
rect 7200 2758 7252 2810
rect 7274 2758 7326 2810
rect 7348 2758 7400 2810
rect 8400 2758 8452 2810
rect 8474 2758 8526 2810
rect 8548 2758 8600 2810
rect 9600 2758 9652 2810
rect 9674 2758 9726 2810
rect 9748 2758 9800 2810
rect 10800 2758 10852 2810
rect 10874 2758 10926 2810
rect 10948 2758 11000 2810
rect 12000 2758 12052 2810
rect 12074 2758 12126 2810
rect 12148 2758 12200 2810
rect 13200 2758 13252 2810
rect 13274 2758 13326 2810
rect 13348 2758 13400 2810
rect 14400 2758 14452 2810
rect 14474 2758 14526 2810
rect 14548 2758 14600 2810
rect 15600 2758 15652 2810
rect 15674 2758 15726 2810
rect 15748 2758 15800 2810
rect 16800 2758 16852 2810
rect 16874 2758 16926 2810
rect 16948 2758 17000 2810
rect 18000 2758 18052 2810
rect 18074 2758 18126 2810
rect 18148 2758 18200 2810
rect 19200 2758 19252 2810
rect 19274 2758 19326 2810
rect 19348 2758 19400 2810
rect 20400 2758 20452 2810
rect 20474 2758 20526 2810
rect 20548 2758 20600 2810
rect 21156 2758 21208 2810
rect 21230 2758 21282 2810
rect 21304 2758 21356 2810
<< metal2 >>
rect 20400 3882 20600 3903
rect 20400 3826 20420 3882
rect 20476 3826 20524 3882
rect 20580 3826 20600 3882
rect 20400 3778 20600 3826
rect 20400 3722 20420 3778
rect 20476 3722 20524 3778
rect 20580 3722 20600 3778
rect 20400 3700 20600 3722
rect 21503 3876 23110 3900
rect 21503 3824 21525 3876
rect 21577 3824 21623 3876
rect 21675 3824 23110 3876
rect 21503 3800 23110 3824
rect 21503 3776 21700 3800
rect 21503 3724 21525 3776
rect 21577 3724 21623 3776
rect 21675 3724 21700 3776
rect 21503 3700 21700 3724
rect 2400 3208 2600 3220
rect 2400 3206 2422 3208
rect 2478 3206 2522 3208
rect 2578 3206 2600 3208
rect 2400 3152 2422 3154
rect 2478 3152 2522 3154
rect 2578 3152 2600 3154
rect 2400 3140 2600 3152
rect 3600 3208 3800 3220
rect 3600 3206 3622 3208
rect 3678 3206 3722 3208
rect 3778 3206 3800 3208
rect 3600 3152 3622 3154
rect 3678 3152 3722 3154
rect 3778 3152 3800 3154
rect 3600 3140 3800 3152
rect 4800 3208 5000 3220
rect 4800 3206 4822 3208
rect 4878 3206 4922 3208
rect 4978 3206 5000 3208
rect 4800 3152 4822 3154
rect 4878 3152 4922 3154
rect 4978 3152 5000 3154
rect 4800 3140 5000 3152
rect 6000 3208 6200 3220
rect 6000 3206 6022 3208
rect 6078 3206 6122 3208
rect 6178 3206 6200 3208
rect 6000 3152 6022 3154
rect 6078 3152 6122 3154
rect 6178 3152 6200 3154
rect 6000 3140 6200 3152
rect 7200 3208 7400 3220
rect 7200 3206 7222 3208
rect 7278 3206 7322 3208
rect 7378 3206 7400 3208
rect 7200 3152 7222 3154
rect 7278 3152 7322 3154
rect 7378 3152 7400 3154
rect 7200 3140 7400 3152
rect 8400 3208 8600 3220
rect 8400 3206 8422 3208
rect 8478 3206 8522 3208
rect 8578 3206 8600 3208
rect 8400 3152 8422 3154
rect 8478 3152 8522 3154
rect 8578 3152 8600 3154
rect 8400 3140 8600 3152
rect 9600 3208 9800 3220
rect 9600 3206 9622 3208
rect 9678 3206 9722 3208
rect 9778 3206 9800 3208
rect 9600 3152 9622 3154
rect 9678 3152 9722 3154
rect 9778 3152 9800 3154
rect 9600 3140 9800 3152
rect 10800 3208 11000 3220
rect 10800 3206 10822 3208
rect 10878 3206 10922 3208
rect 10978 3206 11000 3208
rect 10800 3152 10822 3154
rect 10878 3152 10922 3154
rect 10978 3152 11000 3154
rect 10800 3140 11000 3152
rect 12000 3208 12200 3220
rect 12000 3206 12022 3208
rect 12078 3206 12122 3208
rect 12178 3206 12200 3208
rect 12000 3152 12022 3154
rect 12078 3152 12122 3154
rect 12178 3152 12200 3154
rect 12000 3140 12200 3152
rect 13200 3208 13400 3220
rect 13200 3206 13222 3208
rect 13278 3206 13322 3208
rect 13378 3206 13400 3208
rect 13200 3152 13222 3154
rect 13278 3152 13322 3154
rect 13378 3152 13400 3154
rect 13200 3140 13400 3152
rect 14400 3208 14600 3220
rect 14400 3206 14422 3208
rect 14478 3206 14522 3208
rect 14578 3206 14600 3208
rect 14400 3152 14422 3154
rect 14478 3152 14522 3154
rect 14578 3152 14600 3154
rect 14400 3140 14600 3152
rect 15600 3208 15800 3220
rect 15600 3206 15622 3208
rect 15678 3206 15722 3208
rect 15778 3206 15800 3208
rect 15600 3152 15622 3154
rect 15678 3152 15722 3154
rect 15778 3152 15800 3154
rect 15600 3140 15800 3152
rect 16800 3208 17000 3220
rect 16800 3206 16822 3208
rect 16878 3206 16922 3208
rect 16978 3206 17000 3208
rect 16800 3152 16822 3154
rect 16878 3152 16922 3154
rect 16978 3152 17000 3154
rect 16800 3140 17000 3152
rect 18000 3208 18200 3220
rect 18000 3206 18022 3208
rect 18078 3206 18122 3208
rect 18178 3206 18200 3208
rect 18000 3152 18022 3154
rect 18078 3152 18122 3154
rect 18178 3152 18200 3154
rect 18000 3140 18200 3152
rect 19200 3208 19400 3220
rect 19200 3206 19222 3208
rect 19278 3206 19322 3208
rect 19378 3206 19400 3208
rect 19200 3152 19222 3154
rect 19278 3152 19322 3154
rect 19378 3152 19400 3154
rect 19200 3140 19400 3152
rect 0 2812 200 2824
rect 0 2810 22 2812
rect 78 2810 122 2812
rect 178 2810 200 2812
rect 0 2756 22 2758
rect 78 2756 122 2758
rect 178 2756 200 2758
rect 0 2744 200 2756
rect 1200 2812 1400 2824
rect 1200 2810 1222 2812
rect 1278 2810 1322 2812
rect 1378 2810 1400 2812
rect 1200 2756 1222 2758
rect 1278 2756 1322 2758
rect 1378 2756 1400 2758
rect 1200 2744 1400 2756
rect 2400 2812 2600 2824
rect 2400 2810 2422 2812
rect 2478 2810 2522 2812
rect 2578 2810 2600 2812
rect 2400 2756 2422 2758
rect 2478 2756 2522 2758
rect 2578 2756 2600 2758
rect 2400 2744 2600 2756
rect 3600 2812 3800 2824
rect 3600 2810 3622 2812
rect 3678 2810 3722 2812
rect 3778 2810 3800 2812
rect 3600 2756 3622 2758
rect 3678 2756 3722 2758
rect 3778 2756 3800 2758
rect 3600 2744 3800 2756
rect 4800 2812 5000 2824
rect 4800 2810 4822 2812
rect 4878 2810 4922 2812
rect 4978 2810 5000 2812
rect 4800 2756 4822 2758
rect 4878 2756 4922 2758
rect 4978 2756 5000 2758
rect 4800 2744 5000 2756
rect 6000 2812 6200 2824
rect 6000 2810 6022 2812
rect 6078 2810 6122 2812
rect 6178 2810 6200 2812
rect 6000 2756 6022 2758
rect 6078 2756 6122 2758
rect 6178 2756 6200 2758
rect 6000 2744 6200 2756
rect 7200 2812 7400 2824
rect 7200 2810 7222 2812
rect 7278 2810 7322 2812
rect 7378 2810 7400 2812
rect 7200 2756 7222 2758
rect 7278 2756 7322 2758
rect 7378 2756 7400 2758
rect 7200 2744 7400 2756
rect 8400 2812 8600 2824
rect 8400 2810 8422 2812
rect 8478 2810 8522 2812
rect 8578 2810 8600 2812
rect 8400 2756 8422 2758
rect 8478 2756 8522 2758
rect 8578 2756 8600 2758
rect 8400 2744 8600 2756
rect 9600 2812 9800 2824
rect 9600 2810 9622 2812
rect 9678 2810 9722 2812
rect 9778 2810 9800 2812
rect 9600 2756 9622 2758
rect 9678 2756 9722 2758
rect 9778 2756 9800 2758
rect 9600 2744 9800 2756
rect 10800 2812 11000 2824
rect 10800 2810 10822 2812
rect 10878 2810 10922 2812
rect 10978 2810 11000 2812
rect 10800 2756 10822 2758
rect 10878 2756 10922 2758
rect 10978 2756 11000 2758
rect 10800 2744 11000 2756
rect 12000 2812 12200 2824
rect 12000 2810 12022 2812
rect 12078 2810 12122 2812
rect 12178 2810 12200 2812
rect 12000 2756 12022 2758
rect 12078 2756 12122 2758
rect 12178 2756 12200 2758
rect 12000 2744 12200 2756
rect 13200 2812 13400 2824
rect 13200 2810 13222 2812
rect 13278 2810 13322 2812
rect 13378 2810 13400 2812
rect 13200 2756 13222 2758
rect 13278 2756 13322 2758
rect 13378 2756 13400 2758
rect 13200 2744 13400 2756
rect 14400 2812 14600 2824
rect 14400 2810 14422 2812
rect 14478 2810 14522 2812
rect 14578 2810 14600 2812
rect 14400 2756 14422 2758
rect 14478 2756 14522 2758
rect 14578 2756 14600 2758
rect 14400 2744 14600 2756
rect 15600 2812 15800 2824
rect 15600 2810 15622 2812
rect 15678 2810 15722 2812
rect 15778 2810 15800 2812
rect 15600 2756 15622 2758
rect 15678 2756 15722 2758
rect 15778 2756 15800 2758
rect 15600 2744 15800 2756
rect 16800 2812 17000 2824
rect 16800 2810 16822 2812
rect 16878 2810 16922 2812
rect 16978 2810 17000 2812
rect 16800 2756 16822 2758
rect 16878 2756 16922 2758
rect 16978 2756 17000 2758
rect 16800 2744 17000 2756
rect 18000 2812 18200 2824
rect 18000 2810 18022 2812
rect 18078 2810 18122 2812
rect 18178 2810 18200 2812
rect 18000 2756 18022 2758
rect 18078 2756 18122 2758
rect 18178 2756 18200 2758
rect 18000 2744 18200 2756
rect 19200 2812 19400 2824
rect 19200 2810 19222 2812
rect 19278 2810 19322 2812
rect 19378 2810 19400 2812
rect 19200 2756 19222 2758
rect 19278 2756 19322 2758
rect 19378 2756 19400 2758
rect 19200 2744 19400 2756
rect 20400 2812 20600 2824
rect 20400 2810 20422 2812
rect 20478 2810 20522 2812
rect 20578 2810 20600 2812
rect 20400 2756 20422 2758
rect 20478 2756 20522 2758
rect 20578 2756 20600 2758
rect 20400 2744 20600 2756
rect 21156 2812 21356 2824
rect 21156 2810 21178 2812
rect 21234 2810 21278 2812
rect 21334 2810 21356 2812
rect 21156 2756 21178 2758
rect 21234 2756 21278 2758
rect 21334 2756 21356 2758
rect 21156 2744 21356 2756
<< via2 >>
rect 20420 3880 20476 3882
rect 20420 3828 20422 3880
rect 20422 3828 20474 3880
rect 20474 3828 20476 3880
rect 20420 3826 20476 3828
rect 20524 3880 20580 3882
rect 20524 3828 20526 3880
rect 20526 3828 20578 3880
rect 20578 3828 20580 3880
rect 20524 3826 20580 3828
rect 20420 3776 20476 3778
rect 20420 3724 20422 3776
rect 20422 3724 20474 3776
rect 20474 3724 20476 3776
rect 20420 3722 20476 3724
rect 20524 3776 20580 3778
rect 20524 3724 20526 3776
rect 20526 3724 20578 3776
rect 20578 3724 20580 3776
rect 20524 3722 20580 3724
rect 2422 3206 2478 3208
rect 2522 3206 2578 3208
rect 2422 3154 2452 3206
rect 2452 3154 2474 3206
rect 2474 3154 2478 3206
rect 2522 3154 2526 3206
rect 2526 3154 2548 3206
rect 2548 3154 2578 3206
rect 2422 3152 2478 3154
rect 2522 3152 2578 3154
rect 3622 3206 3678 3208
rect 3722 3206 3778 3208
rect 3622 3154 3652 3206
rect 3652 3154 3674 3206
rect 3674 3154 3678 3206
rect 3722 3154 3726 3206
rect 3726 3154 3748 3206
rect 3748 3154 3778 3206
rect 3622 3152 3678 3154
rect 3722 3152 3778 3154
rect 4822 3206 4878 3208
rect 4922 3206 4978 3208
rect 4822 3154 4852 3206
rect 4852 3154 4874 3206
rect 4874 3154 4878 3206
rect 4922 3154 4926 3206
rect 4926 3154 4948 3206
rect 4948 3154 4978 3206
rect 4822 3152 4878 3154
rect 4922 3152 4978 3154
rect 6022 3206 6078 3208
rect 6122 3206 6178 3208
rect 6022 3154 6052 3206
rect 6052 3154 6074 3206
rect 6074 3154 6078 3206
rect 6122 3154 6126 3206
rect 6126 3154 6148 3206
rect 6148 3154 6178 3206
rect 6022 3152 6078 3154
rect 6122 3152 6178 3154
rect 7222 3206 7278 3208
rect 7322 3206 7378 3208
rect 7222 3154 7252 3206
rect 7252 3154 7274 3206
rect 7274 3154 7278 3206
rect 7322 3154 7326 3206
rect 7326 3154 7348 3206
rect 7348 3154 7378 3206
rect 7222 3152 7278 3154
rect 7322 3152 7378 3154
rect 8422 3206 8478 3208
rect 8522 3206 8578 3208
rect 8422 3154 8452 3206
rect 8452 3154 8474 3206
rect 8474 3154 8478 3206
rect 8522 3154 8526 3206
rect 8526 3154 8548 3206
rect 8548 3154 8578 3206
rect 8422 3152 8478 3154
rect 8522 3152 8578 3154
rect 9622 3206 9678 3208
rect 9722 3206 9778 3208
rect 9622 3154 9652 3206
rect 9652 3154 9674 3206
rect 9674 3154 9678 3206
rect 9722 3154 9726 3206
rect 9726 3154 9748 3206
rect 9748 3154 9778 3206
rect 9622 3152 9678 3154
rect 9722 3152 9778 3154
rect 10822 3206 10878 3208
rect 10922 3206 10978 3208
rect 10822 3154 10852 3206
rect 10852 3154 10874 3206
rect 10874 3154 10878 3206
rect 10922 3154 10926 3206
rect 10926 3154 10948 3206
rect 10948 3154 10978 3206
rect 10822 3152 10878 3154
rect 10922 3152 10978 3154
rect 12022 3206 12078 3208
rect 12122 3206 12178 3208
rect 12022 3154 12052 3206
rect 12052 3154 12074 3206
rect 12074 3154 12078 3206
rect 12122 3154 12126 3206
rect 12126 3154 12148 3206
rect 12148 3154 12178 3206
rect 12022 3152 12078 3154
rect 12122 3152 12178 3154
rect 13222 3206 13278 3208
rect 13322 3206 13378 3208
rect 13222 3154 13252 3206
rect 13252 3154 13274 3206
rect 13274 3154 13278 3206
rect 13322 3154 13326 3206
rect 13326 3154 13348 3206
rect 13348 3154 13378 3206
rect 13222 3152 13278 3154
rect 13322 3152 13378 3154
rect 14422 3206 14478 3208
rect 14522 3206 14578 3208
rect 14422 3154 14452 3206
rect 14452 3154 14474 3206
rect 14474 3154 14478 3206
rect 14522 3154 14526 3206
rect 14526 3154 14548 3206
rect 14548 3154 14578 3206
rect 14422 3152 14478 3154
rect 14522 3152 14578 3154
rect 15622 3206 15678 3208
rect 15722 3206 15778 3208
rect 15622 3154 15652 3206
rect 15652 3154 15674 3206
rect 15674 3154 15678 3206
rect 15722 3154 15726 3206
rect 15726 3154 15748 3206
rect 15748 3154 15778 3206
rect 15622 3152 15678 3154
rect 15722 3152 15778 3154
rect 16822 3206 16878 3208
rect 16922 3206 16978 3208
rect 16822 3154 16852 3206
rect 16852 3154 16874 3206
rect 16874 3154 16878 3206
rect 16922 3154 16926 3206
rect 16926 3154 16948 3206
rect 16948 3154 16978 3206
rect 16822 3152 16878 3154
rect 16922 3152 16978 3154
rect 18022 3206 18078 3208
rect 18122 3206 18178 3208
rect 18022 3154 18052 3206
rect 18052 3154 18074 3206
rect 18074 3154 18078 3206
rect 18122 3154 18126 3206
rect 18126 3154 18148 3206
rect 18148 3154 18178 3206
rect 18022 3152 18078 3154
rect 18122 3152 18178 3154
rect 19222 3206 19278 3208
rect 19322 3206 19378 3208
rect 19222 3154 19252 3206
rect 19252 3154 19274 3206
rect 19274 3154 19278 3206
rect 19322 3154 19326 3206
rect 19326 3154 19348 3206
rect 19348 3154 19378 3206
rect 19222 3152 19278 3154
rect 19322 3152 19378 3154
rect 22 2810 78 2812
rect 122 2810 178 2812
rect 22 2758 52 2810
rect 52 2758 74 2810
rect 74 2758 78 2810
rect 122 2758 126 2810
rect 126 2758 148 2810
rect 148 2758 178 2810
rect 22 2756 78 2758
rect 122 2756 178 2758
rect 1222 2810 1278 2812
rect 1322 2810 1378 2812
rect 1222 2758 1252 2810
rect 1252 2758 1274 2810
rect 1274 2758 1278 2810
rect 1322 2758 1326 2810
rect 1326 2758 1348 2810
rect 1348 2758 1378 2810
rect 1222 2756 1278 2758
rect 1322 2756 1378 2758
rect 2422 2810 2478 2812
rect 2522 2810 2578 2812
rect 2422 2758 2452 2810
rect 2452 2758 2474 2810
rect 2474 2758 2478 2810
rect 2522 2758 2526 2810
rect 2526 2758 2548 2810
rect 2548 2758 2578 2810
rect 2422 2756 2478 2758
rect 2522 2756 2578 2758
rect 3622 2810 3678 2812
rect 3722 2810 3778 2812
rect 3622 2758 3652 2810
rect 3652 2758 3674 2810
rect 3674 2758 3678 2810
rect 3722 2758 3726 2810
rect 3726 2758 3748 2810
rect 3748 2758 3778 2810
rect 3622 2756 3678 2758
rect 3722 2756 3778 2758
rect 4822 2810 4878 2812
rect 4922 2810 4978 2812
rect 4822 2758 4852 2810
rect 4852 2758 4874 2810
rect 4874 2758 4878 2810
rect 4922 2758 4926 2810
rect 4926 2758 4948 2810
rect 4948 2758 4978 2810
rect 4822 2756 4878 2758
rect 4922 2756 4978 2758
rect 6022 2810 6078 2812
rect 6122 2810 6178 2812
rect 6022 2758 6052 2810
rect 6052 2758 6074 2810
rect 6074 2758 6078 2810
rect 6122 2758 6126 2810
rect 6126 2758 6148 2810
rect 6148 2758 6178 2810
rect 6022 2756 6078 2758
rect 6122 2756 6178 2758
rect 7222 2810 7278 2812
rect 7322 2810 7378 2812
rect 7222 2758 7252 2810
rect 7252 2758 7274 2810
rect 7274 2758 7278 2810
rect 7322 2758 7326 2810
rect 7326 2758 7348 2810
rect 7348 2758 7378 2810
rect 7222 2756 7278 2758
rect 7322 2756 7378 2758
rect 8422 2810 8478 2812
rect 8522 2810 8578 2812
rect 8422 2758 8452 2810
rect 8452 2758 8474 2810
rect 8474 2758 8478 2810
rect 8522 2758 8526 2810
rect 8526 2758 8548 2810
rect 8548 2758 8578 2810
rect 8422 2756 8478 2758
rect 8522 2756 8578 2758
rect 9622 2810 9678 2812
rect 9722 2810 9778 2812
rect 9622 2758 9652 2810
rect 9652 2758 9674 2810
rect 9674 2758 9678 2810
rect 9722 2758 9726 2810
rect 9726 2758 9748 2810
rect 9748 2758 9778 2810
rect 9622 2756 9678 2758
rect 9722 2756 9778 2758
rect 10822 2810 10878 2812
rect 10922 2810 10978 2812
rect 10822 2758 10852 2810
rect 10852 2758 10874 2810
rect 10874 2758 10878 2810
rect 10922 2758 10926 2810
rect 10926 2758 10948 2810
rect 10948 2758 10978 2810
rect 10822 2756 10878 2758
rect 10922 2756 10978 2758
rect 12022 2810 12078 2812
rect 12122 2810 12178 2812
rect 12022 2758 12052 2810
rect 12052 2758 12074 2810
rect 12074 2758 12078 2810
rect 12122 2758 12126 2810
rect 12126 2758 12148 2810
rect 12148 2758 12178 2810
rect 12022 2756 12078 2758
rect 12122 2756 12178 2758
rect 13222 2810 13278 2812
rect 13322 2810 13378 2812
rect 13222 2758 13252 2810
rect 13252 2758 13274 2810
rect 13274 2758 13278 2810
rect 13322 2758 13326 2810
rect 13326 2758 13348 2810
rect 13348 2758 13378 2810
rect 13222 2756 13278 2758
rect 13322 2756 13378 2758
rect 14422 2810 14478 2812
rect 14522 2810 14578 2812
rect 14422 2758 14452 2810
rect 14452 2758 14474 2810
rect 14474 2758 14478 2810
rect 14522 2758 14526 2810
rect 14526 2758 14548 2810
rect 14548 2758 14578 2810
rect 14422 2756 14478 2758
rect 14522 2756 14578 2758
rect 15622 2810 15678 2812
rect 15722 2810 15778 2812
rect 15622 2758 15652 2810
rect 15652 2758 15674 2810
rect 15674 2758 15678 2810
rect 15722 2758 15726 2810
rect 15726 2758 15748 2810
rect 15748 2758 15778 2810
rect 15622 2756 15678 2758
rect 15722 2756 15778 2758
rect 16822 2810 16878 2812
rect 16922 2810 16978 2812
rect 16822 2758 16852 2810
rect 16852 2758 16874 2810
rect 16874 2758 16878 2810
rect 16922 2758 16926 2810
rect 16926 2758 16948 2810
rect 16948 2758 16978 2810
rect 16822 2756 16878 2758
rect 16922 2756 16978 2758
rect 18022 2810 18078 2812
rect 18122 2810 18178 2812
rect 18022 2758 18052 2810
rect 18052 2758 18074 2810
rect 18074 2758 18078 2810
rect 18122 2758 18126 2810
rect 18126 2758 18148 2810
rect 18148 2758 18178 2810
rect 18022 2756 18078 2758
rect 18122 2756 18178 2758
rect 19222 2810 19278 2812
rect 19322 2810 19378 2812
rect 19222 2758 19252 2810
rect 19252 2758 19274 2810
rect 19274 2758 19278 2810
rect 19322 2758 19326 2810
rect 19326 2758 19348 2810
rect 19348 2758 19378 2810
rect 19222 2756 19278 2758
rect 19322 2756 19378 2758
rect 20422 2810 20478 2812
rect 20522 2810 20578 2812
rect 20422 2758 20452 2810
rect 20452 2758 20474 2810
rect 20474 2758 20478 2810
rect 20522 2758 20526 2810
rect 20526 2758 20548 2810
rect 20548 2758 20578 2810
rect 20422 2756 20478 2758
rect 20522 2756 20578 2758
rect 21178 2810 21234 2812
rect 21278 2810 21334 2812
rect 21178 2758 21208 2810
rect 21208 2758 21230 2810
rect 21230 2758 21234 2810
rect 21278 2758 21282 2810
rect 21282 2758 21304 2810
rect 21304 2758 21334 2810
rect 21178 2756 21234 2758
rect 21278 2756 21334 2758
<< metal3 >>
rect 20400 3882 20600 3903
rect 20400 3826 20420 3882
rect 20476 3826 20524 3882
rect 20580 3826 20600 3882
rect 20400 3778 20600 3826
rect 20400 3722 20420 3778
rect 20476 3722 20524 3778
rect 20580 3722 20600 3778
rect 2400 3208 2600 3230
rect 2400 3152 2422 3208
rect 2478 3152 2522 3208
rect 2578 3152 2600 3208
rect 2400 3134 2600 3152
rect 3600 3208 3800 3230
rect 3600 3152 3622 3208
rect 3678 3152 3722 3208
rect 3778 3152 3800 3208
rect 3600 3134 3800 3152
rect 4800 3208 5000 3230
rect 4800 3152 4822 3208
rect 4878 3152 4922 3208
rect 4978 3152 5000 3208
rect 4800 3134 5000 3152
rect 6000 3208 6200 3230
rect 6000 3152 6022 3208
rect 6078 3152 6122 3208
rect 6178 3152 6200 3208
rect 6000 3134 6200 3152
rect 7200 3208 7400 3230
rect 7200 3152 7222 3208
rect 7278 3152 7322 3208
rect 7378 3152 7400 3208
rect 7200 3134 7400 3152
rect 8400 3208 8600 3230
rect 8400 3152 8422 3208
rect 8478 3152 8522 3208
rect 8578 3152 8600 3208
rect 8400 3134 8600 3152
rect 9600 3208 9800 3230
rect 9600 3152 9622 3208
rect 9678 3152 9722 3208
rect 9778 3152 9800 3208
rect 9600 3134 9800 3152
rect 10800 3208 11000 3230
rect 10800 3152 10822 3208
rect 10878 3152 10922 3208
rect 10978 3152 11000 3208
rect 10800 3134 11000 3152
rect 12000 3208 12200 3230
rect 12000 3152 12022 3208
rect 12078 3152 12122 3208
rect 12178 3152 12200 3208
rect 12000 3134 12200 3152
rect 13200 3208 13400 3230
rect 13200 3152 13222 3208
rect 13278 3152 13322 3208
rect 13378 3152 13400 3208
rect 13200 3134 13400 3152
rect 14400 3208 14600 3230
rect 14400 3152 14422 3208
rect 14478 3152 14522 3208
rect 14578 3152 14600 3208
rect 14400 3134 14600 3152
rect 15600 3208 15800 3230
rect 15600 3152 15622 3208
rect 15678 3152 15722 3208
rect 15778 3152 15800 3208
rect 15600 3134 15800 3152
rect 16800 3208 17000 3230
rect 16800 3152 16822 3208
rect 16878 3152 16922 3208
rect 16978 3152 17000 3208
rect 16800 3134 17000 3152
rect 18000 3208 18200 3230
rect 18000 3152 18022 3208
rect 18078 3152 18122 3208
rect 18178 3152 18200 3208
rect 18000 3134 18200 3152
rect 19200 3208 19400 3230
rect 19200 3152 19222 3208
rect 19278 3152 19322 3208
rect 19378 3152 19400 3208
rect 19200 3134 19400 3152
rect 20400 3134 20600 3722
rect 0 2834 21356 3134
rect 0 2812 200 2834
rect 0 2756 22 2812
rect 78 2756 122 2812
rect 178 2756 200 2812
rect 0 2738 200 2756
rect 1200 2812 1400 2834
rect 1200 2756 1222 2812
rect 1278 2756 1322 2812
rect 1378 2756 1400 2812
rect 1200 2738 1400 2756
rect 2400 2812 2600 2834
rect 2400 2756 2422 2812
rect 2478 2756 2522 2812
rect 2578 2756 2600 2812
rect 2400 2738 2600 2756
rect 3600 2812 3800 2834
rect 3600 2756 3622 2812
rect 3678 2756 3722 2812
rect 3778 2756 3800 2812
rect 3600 2738 3800 2756
rect 4800 2812 5000 2834
rect 4800 2756 4822 2812
rect 4878 2756 4922 2812
rect 4978 2756 5000 2812
rect 4800 2738 5000 2756
rect 6000 2812 6200 2834
rect 6000 2756 6022 2812
rect 6078 2756 6122 2812
rect 6178 2756 6200 2812
rect 6000 2738 6200 2756
rect 7200 2812 7400 2834
rect 7200 2756 7222 2812
rect 7278 2756 7322 2812
rect 7378 2756 7400 2812
rect 7200 2738 7400 2756
rect 8400 2812 8600 2834
rect 8400 2756 8422 2812
rect 8478 2756 8522 2812
rect 8578 2756 8600 2812
rect 8400 2738 8600 2756
rect 9600 2812 9800 2834
rect 9600 2756 9622 2812
rect 9678 2756 9722 2812
rect 9778 2756 9800 2812
rect 9600 2738 9800 2756
rect 10800 2812 11000 2834
rect 10800 2756 10822 2812
rect 10878 2756 10922 2812
rect 10978 2756 11000 2812
rect 10800 2738 11000 2756
rect 12000 2812 12200 2834
rect 12000 2756 12022 2812
rect 12078 2756 12122 2812
rect 12178 2756 12200 2812
rect 12000 2738 12200 2756
rect 13200 2812 13400 2834
rect 13200 2756 13222 2812
rect 13278 2756 13322 2812
rect 13378 2756 13400 2812
rect 13200 2738 13400 2756
rect 14400 2812 14600 2834
rect 14400 2756 14422 2812
rect 14478 2756 14522 2812
rect 14578 2756 14600 2812
rect 14400 2738 14600 2756
rect 15600 2812 15800 2834
rect 15600 2756 15622 2812
rect 15678 2756 15722 2812
rect 15778 2756 15800 2812
rect 15600 2738 15800 2756
rect 16800 2812 17000 2834
rect 16800 2756 16822 2812
rect 16878 2756 16922 2812
rect 16978 2756 17000 2812
rect 16800 2738 17000 2756
rect 18000 2812 18200 2834
rect 18000 2756 18022 2812
rect 18078 2756 18122 2812
rect 18178 2756 18200 2812
rect 18000 2738 18200 2756
rect 19200 2812 19400 2834
rect 19200 2756 19222 2812
rect 19278 2756 19322 2812
rect 19378 2756 19400 2812
rect 19200 2738 19400 2756
rect 20400 2812 20600 2834
rect 20400 2756 20422 2812
rect 20478 2756 20522 2812
rect 20578 2756 20600 2812
rect 20400 2738 20600 2756
rect 21156 2812 21356 2834
rect 21156 2756 21178 2812
rect 21234 2756 21278 2812
rect 21334 2756 21356 2812
rect 21156 2738 21356 2756
use inv  inv_0
timestamp 1623637110
transform -1 0 3246 0 -1 4834
box -400 1960 3246 4834
use inv  inv_2
timestamp 1623637110
transform -1 0 6788 0 -1 4834
box -400 1960 3246 4834
use inv  inv_1
timestamp 1623637110
transform -1 0 10330 0 -1 4834
box -400 1960 3246 4834
use inv  inv_3
timestamp 1623637110
transform -1 0 13872 0 -1 4834
box -400 1960 3246 4834
use inv  inv_4
timestamp 1623637110
transform -1 0 17414 0 -1 4834
box -400 1960 3246 4834
use inv  inv_5
timestamp 1623637110
transform -1 0 20956 0 -1 4834
box -400 1960 3246 4834
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1630125002
transform 1 0 -162 0 1 4560
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1630125002
transform 1 0 637 0 1 4560
box -38 -48 314 592
use inv  inv_6
timestamp 1623637110
transform 1 0 2096 0 1 1134
box -400 1960 3246 4834
use inv  inv_7
timestamp 1623637110
transform 1 0 5638 0 1 1134
box -400 1960 3246 4834
use inv  inv_8
timestamp 1623637110
transform 1 0 9180 0 1 1134
box -400 1960 3246 4834
use inv  inv_9
timestamp 1623637110
transform 1 0 12722 0 1 1134
box -400 1960 3246 4834
use inv  inv_10
timestamp 1623637110
transform 1 0 16264 0 1 1134
box -400 1960 3246 4834
use res_poly  res_poly_0
timestamp 1637941551
transform 1 0 20200 0 1 3900
box 0 -6 400 976
use res_poly  res_poly_1
timestamp 1637941551
transform 0 1 20600 -1 0 3900
box 0 -6 400 976
<< labels >>
flabel metal1 s 5254 4790 5326 4862 1 FreeSans 250 0 0 0 p[6]
port 1 nsew
flabel metal1 s 19510 4790 19582 4862 1 FreeSans 250 0 0 0 p[10]
port 2 nsew
flabel metal1 s 17728 1650 17800 1722 1 FreeSans 250 0 0 0 pn[0]
port 3 nsew
flabel metal1 s 14182 1650 14254 1722 1 FreeSans 250 0 0 0 pn[1]
port 4 nsew
flabel metal1 s 10634 1650 10706 1722 1 FreeSans 250 0 0 0 pn[2]
port 5 nsew
flabel metal1 s 7104 1650 7176 1722 1 FreeSans 250 0 0 0 pn[3]
port 6 nsew
flabel metal1 s 3554 1650 3626 1722 1 FreeSans 250 0 0 0 pn[4]
port 7 nsew
flabel metal1 s -72 1650 0 1722 1 FreeSans 250 0 0 0 pn[5]
port 8 nsew
flabel metal1 s 5254 4246 5326 4318 1 FreeSans 250 0 0 0 pn[6]
port 9 nsew
flabel metal1 s 8798 4246 8870 4318 1 FreeSans 250 0 0 0 pn[7]
port 10 nsew
flabel metal1 s 12334 4246 12406 4318 1 FreeSans 250 0 0 0 pn[8]
port 11 nsew
flabel metal1 s 15878 4246 15950 4318 1 FreeSans 250 0 0 0 pn[9]
port 12 nsew
flabel metal1 s 19510 4246 19582 4318 1 FreeSans 250 0 0 0 pn[10]
port 13 nsew
flabel metal2 s 21600 3800 21700 3900 1 FreeSans 250 0 0 0 input_analog
port 14 nsew
flabel metal3 s 20400 3498 20502 3600 1 FreeSans 250 0 0 0 v_ctr
port 15 nsew
flabel metal1 s -200 4512 -104 4608 1 FreeSans 250 0 0 0 vssd2
port 16 nsew
flabel metal1 s -200 5056 -104 5152 1 FreeSans 250 0 0 0 vccd2
port 17 nsew
flabel metal1 s 1680 5854 1776 5950 1 FreeSans 250 0 0 0 vccd2
port 17 nsew
flabel metal1 s 20524 4804 20596 4876 1 FreeSans 250 0 0 0 vssd2
port 16 nsew
flabel metal1 s 10650 1106 10722 1178 1 FreeSans 250 0 0 0 p[2]        
port 18 nsew
flabel metal1 s 14182 1106 14254 1178 1 FreeSans 250 0 0 0 p[1]        
port 19 nsew
flabel metal1 s 15878 4790 15950 4862 1 FreeSans 250 0 0 0 p[9]
port 20 nsew
flabel metal1 s 12334 4790 12406 4862 1 FreeSans 250 0 0 0 p[8]
port 21 nsew
<< end >>
