magic
tech sky130A
timestamp 1623055983
<< pwell >>
rect -98 -105 288 605
<< nmos >>
rect 0 0 190 500
<< ndiff >>
rect -29 482 0 500
rect -29 462 -23 482
rect -6 462 0 482
rect -29 445 0 462
rect -29 425 -23 445
rect -6 425 0 445
rect -29 408 0 425
rect -29 388 -23 408
rect -6 388 0 408
rect -29 371 0 388
rect -29 351 -23 371
rect -6 351 0 371
rect -29 334 0 351
rect -29 314 -23 334
rect -6 314 0 334
rect -29 297 0 314
rect -29 277 -23 297
rect -6 277 0 297
rect -29 260 0 277
rect -29 240 -23 260
rect -6 240 0 260
rect -29 222 0 240
rect -29 202 -23 222
rect -6 202 0 222
rect -29 185 0 202
rect -29 165 -23 185
rect -6 165 0 185
rect -29 148 0 165
rect -29 128 -23 148
rect -6 128 0 148
rect -29 111 0 128
rect -29 91 -23 111
rect -6 91 0 111
rect -29 74 0 91
rect -29 54 -23 74
rect -6 54 0 74
rect -29 37 0 54
rect -29 17 -23 37
rect -6 17 0 37
rect -29 0 0 17
rect 190 482 219 500
rect 190 462 196 482
rect 213 462 219 482
rect 190 445 219 462
rect 190 425 196 445
rect 213 425 219 445
rect 190 408 219 425
rect 190 388 196 408
rect 213 388 219 408
rect 190 371 219 388
rect 190 351 196 371
rect 213 351 219 371
rect 190 334 219 351
rect 190 314 196 334
rect 213 314 219 334
rect 190 297 219 314
rect 190 277 196 297
rect 213 277 219 297
rect 190 260 219 277
rect 190 240 196 260
rect 213 240 219 260
rect 190 222 219 240
rect 190 202 196 222
rect 213 202 219 222
rect 190 185 219 202
rect 190 165 196 185
rect 213 165 219 185
rect 190 148 219 165
rect 190 128 196 148
rect 213 128 219 148
rect 190 111 219 128
rect 190 91 196 111
rect 213 91 219 111
rect 190 74 219 91
rect 190 54 196 74
rect 213 54 219 74
rect 190 37 219 54
rect 190 17 196 37
rect 213 17 219 37
rect 190 0 219 17
<< ndiffc >>
rect -23 462 -6 482
rect -23 425 -6 445
rect -23 388 -6 408
rect -23 351 -6 371
rect -23 314 -6 334
rect -23 277 -6 297
rect -23 240 -6 260
rect -23 202 -6 222
rect -23 165 -6 185
rect -23 128 -6 148
rect -23 91 -6 111
rect -23 54 -6 74
rect -23 17 -6 37
rect 196 462 213 482
rect 196 425 213 445
rect 196 388 213 408
rect 196 351 213 371
rect 196 314 213 334
rect 196 277 213 297
rect 196 240 213 260
rect 196 202 213 222
rect 196 165 213 185
rect 196 128 213 148
rect 196 91 213 111
rect 196 54 213 74
rect 196 17 213 37
<< poly >>
rect 0 500 190 544
rect 0 -13 190 0
<< locali >>
rect -23 482 -6 502
rect -23 445 -6 462
rect -23 408 -6 425
rect -23 371 -6 388
rect -23 334 -6 351
rect -23 297 -6 314
rect -23 260 -6 277
rect -23 222 -6 240
rect -23 185 -6 202
rect -23 148 -6 165
rect -23 111 -6 128
rect -23 74 -6 91
rect -23 37 -6 54
rect -23 -2 -6 17
rect 196 482 213 502
rect 196 445 213 462
rect 196 408 213 425
rect 196 371 213 388
rect 196 334 213 351
rect 196 297 213 314
rect 196 260 213 277
rect 196 222 213 240
rect 196 185 213 202
rect 196 148 213 165
rect 196 111 213 128
rect 196 74 213 91
rect 196 37 213 54
rect 196 -2 213 17
<< end >>
