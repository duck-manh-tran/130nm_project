magic
tech sky130A
magscale 1 2
timestamp 1637580353
<< nwell >>
rect 19820 4234 19836 4420
<< pwell >>
rect 528 3668 1752 3700
rect 18924 3668 21196 3700
rect 528 3332 21196 3668
<< pdiff >>
rect 19848 4526 20018 4602
rect 19860 4502 20018 4526
rect 19860 4466 19882 4502
rect 19918 4466 20018 4502
rect 19860 4445 20018 4466
rect 19942 4432 20018 4445
<< pdiffc >>
rect 19882 4466 19918 4502
<< psubdiff >>
rect 4618 7100 4640 7160
rect 4700 7100 4760 7160
rect 4820 7100 4880 7160
rect 4940 7100 5000 7160
rect 5060 7100 5082 7160
rect 10144 7100 10160 7160
rect 10220 7100 10236 7160
rect 10384 7100 10400 7160
rect 10460 7100 10476 7160
rect 10504 7100 10520 7160
rect 10580 7100 10596 7160
rect 15778 7100 15800 7160
rect 15860 7100 15920 7160
rect 15980 7100 16040 7160
rect 16100 7100 16160 7160
rect 16220 7100 16242 7160
rect 4598 -160 4620 -100
rect 4680 -160 4740 -100
rect 4800 -160 4860 -100
rect 4920 -160 4980 -100
rect 5040 -160 5062 -100
rect 10118 -160 10140 -100
rect 10200 -160 10260 -100
rect 10320 -160 10380 -100
rect 10440 -160 10500 -100
rect 10560 -160 10582 -100
rect 15758 -160 15780 -100
rect 15840 -160 15900 -100
rect 15960 -160 16020 -100
rect 16080 -160 16140 -100
rect 16200 -160 16222 -100
<< psubdiffcont >>
rect 4640 7100 4700 7160
rect 4760 7100 4820 7160
rect 4880 7100 4940 7160
rect 5000 7100 5060 7160
rect 10160 7100 10220 7160
rect 10400 7100 10460 7160
rect 10520 7100 10580 7160
rect 15800 7100 15860 7160
rect 15920 7100 15980 7160
rect 16040 7100 16100 7160
rect 16160 7100 16220 7160
rect 4620 -160 4680 -100
rect 4740 -160 4800 -100
rect 4860 -160 4920 -100
rect 4980 -160 5040 -100
rect 10140 -160 10200 -100
rect 10260 -160 10320 -100
rect 10380 -160 10440 -100
rect 10500 -160 10560 -100
rect 15780 -160 15840 -100
rect 15900 -160 15960 -100
rect 16020 -160 16080 -100
rect 16140 -160 16200 -100
<< locali >>
rect 4618 7100 4636 7160
rect 4704 7100 4756 7160
rect 4824 7100 4876 7160
rect 4944 7100 4996 7160
rect 5064 7100 5082 7160
rect 10144 7100 10156 7160
rect 10224 7100 10236 7160
rect 10384 7100 10396 7160
rect 10464 7100 10476 7160
rect 10504 7100 10516 7160
rect 10584 7100 10596 7160
rect 15778 7100 15796 7160
rect 15864 7100 15916 7160
rect 15984 7100 16036 7160
rect 16104 7100 16156 7160
rect 16224 7100 16242 7160
rect 19848 4526 20018 4602
rect 19860 4504 20018 4526
rect 19860 4464 19880 4504
rect 19920 4464 20018 4504
rect 19860 4445 20018 4464
rect 19942 4432 20018 4445
rect 4598 -160 4616 -100
rect 4684 -160 4736 -100
rect 4804 -160 4856 -100
rect 4924 -160 4976 -100
rect 5044 -160 5062 -100
rect 10118 -160 10136 -100
rect 10204 -160 10256 -100
rect 10324 -160 10376 -100
rect 10444 -160 10496 -100
rect 10564 -160 10582 -100
rect 15758 -160 15776 -100
rect 15844 -160 15896 -100
rect 15964 -160 16016 -100
rect 16084 -160 16136 -100
rect 16204 -160 16222 -100
<< viali >>
rect 4636 7160 4704 7164
rect 4756 7160 4824 7164
rect 4876 7160 4944 7164
rect 4996 7160 5064 7164
rect 10156 7160 10224 7164
rect 4636 7100 4640 7160
rect 4640 7100 4700 7160
rect 4700 7100 4704 7160
rect 4756 7100 4760 7160
rect 4760 7100 4820 7160
rect 4820 7100 4824 7160
rect 4876 7100 4880 7160
rect 4880 7100 4940 7160
rect 4940 7100 4944 7160
rect 4996 7100 5000 7160
rect 5000 7100 5060 7160
rect 5060 7100 5064 7160
rect 10156 7100 10160 7160
rect 10160 7100 10220 7160
rect 10220 7100 10224 7160
rect 4636 7096 4704 7100
rect 4756 7096 4824 7100
rect 4876 7096 4944 7100
rect 4996 7096 5064 7100
rect 10156 7096 10224 7100
rect 10276 7096 10344 7164
rect 10396 7160 10464 7164
rect 10516 7160 10584 7164
rect 15796 7160 15864 7164
rect 15916 7160 15984 7164
rect 16036 7160 16104 7164
rect 16156 7160 16224 7164
rect 10396 7100 10400 7160
rect 10400 7100 10460 7160
rect 10460 7100 10464 7160
rect 10516 7100 10520 7160
rect 10520 7100 10580 7160
rect 10580 7100 10584 7160
rect 15796 7100 15800 7160
rect 15800 7100 15860 7160
rect 15860 7100 15864 7160
rect 15916 7100 15920 7160
rect 15920 7100 15980 7160
rect 15980 7100 15984 7160
rect 16036 7100 16040 7160
rect 16040 7100 16100 7160
rect 16100 7100 16104 7160
rect 16156 7100 16160 7160
rect 16160 7100 16220 7160
rect 16220 7100 16224 7160
rect 10396 7096 10464 7100
rect 10516 7096 10584 7100
rect 15796 7096 15864 7100
rect 15916 7096 15984 7100
rect 16036 7096 16104 7100
rect 16156 7096 16224 7100
rect 19880 4502 19920 4504
rect 19880 4466 19882 4502
rect 19882 4466 19918 4502
rect 19918 4466 19920 4502
rect 19880 4464 19920 4466
rect 4616 -100 4684 -96
rect 4736 -100 4804 -96
rect 4856 -100 4924 -96
rect 4976 -100 5044 -96
rect 10136 -100 10204 -96
rect 10256 -100 10324 -96
rect 10376 -100 10444 -96
rect 10496 -100 10564 -96
rect 15776 -100 15844 -96
rect 15896 -100 15964 -96
rect 16016 -100 16084 -96
rect 16136 -100 16204 -96
rect 4616 -160 4620 -100
rect 4620 -160 4680 -100
rect 4680 -160 4684 -100
rect 4736 -160 4740 -100
rect 4740 -160 4800 -100
rect 4800 -160 4804 -100
rect 4856 -160 4860 -100
rect 4860 -160 4920 -100
rect 4920 -160 4924 -100
rect 4976 -160 4980 -100
rect 4980 -160 5040 -100
rect 5040 -160 5044 -100
rect 10136 -160 10140 -100
rect 10140 -160 10200 -100
rect 10200 -160 10204 -100
rect 10256 -160 10260 -100
rect 10260 -160 10320 -100
rect 10320 -160 10324 -100
rect 10376 -160 10380 -100
rect 10380 -160 10440 -100
rect 10440 -160 10444 -100
rect 10496 -160 10500 -100
rect 10500 -160 10560 -100
rect 10560 -160 10564 -100
rect 15776 -160 15780 -100
rect 15780 -160 15840 -100
rect 15840 -160 15844 -100
rect 15896 -160 15900 -100
rect 15900 -160 15960 -100
rect 15960 -160 15964 -100
rect 16016 -160 16020 -100
rect 16020 -160 16080 -100
rect 16080 -160 16084 -100
rect 16136 -160 16140 -100
rect 16140 -160 16200 -100
rect 16200 -160 16204 -100
rect 4616 -164 4684 -160
rect 4736 -164 4804 -160
rect 4856 -164 4924 -160
rect 4976 -164 5044 -160
rect 10136 -164 10204 -160
rect 10256 -164 10324 -160
rect 10376 -164 10444 -160
rect 10496 -164 10564 -160
rect 15776 -164 15844 -160
rect 15896 -164 15964 -160
rect 16016 -164 16084 -160
rect 16136 -164 16204 -160
<< metal1 >>
rect 4618 7168 5082 7180
rect 4618 7092 4632 7168
rect 4708 7092 4752 7168
rect 4828 7092 4872 7168
rect 4948 7092 4992 7168
rect 5068 7092 5082 7168
rect 4618 7080 5082 7092
rect 10138 7168 10602 7180
rect 10138 7092 10152 7168
rect 10228 7092 10272 7168
rect 10348 7092 10392 7168
rect 10468 7092 10512 7168
rect 10588 7092 10602 7168
rect 10138 7080 10602 7092
rect 15778 7168 16242 7180
rect 15778 7092 15792 7168
rect 15868 7092 15912 7168
rect 15988 7092 16032 7168
rect 16108 7092 16152 7168
rect 16228 7092 16242 7168
rect 15778 7080 16242 7092
rect 18914 6924 19000 6938
rect 7422 6918 7498 6924
rect 7422 6854 7428 6918
rect 7492 6854 7498 6918
rect 7422 6848 7498 6854
rect 7566 6918 7642 6924
rect 7566 6854 7572 6918
rect 7636 6854 7642 6918
rect 7566 6848 7642 6854
rect 7710 6918 7786 6924
rect 7710 6854 7716 6918
rect 7780 6854 7786 6918
rect 7710 6848 7786 6854
rect 12946 6918 13022 6924
rect 12946 6854 12952 6918
rect 13016 6854 13022 6918
rect 12946 6848 13022 6854
rect 13090 6918 13166 6924
rect 13090 6854 13096 6918
rect 13160 6854 13166 6918
rect 13090 6848 13166 6854
rect 13250 6918 13326 6924
rect 13250 6854 13256 6918
rect 13320 6854 13326 6918
rect 13250 6848 13326 6854
rect 18558 6918 18634 6924
rect 18558 6854 18564 6918
rect 18628 6854 18634 6918
rect 18558 6848 18634 6854
rect 18702 6918 18778 6924
rect 18702 6854 18708 6918
rect 18772 6854 18778 6918
rect 18702 6848 18778 6854
rect 18842 6918 19000 6924
rect 18842 6854 18848 6918
rect 18912 6854 19000 6918
rect 18842 6848 19000 6854
rect 18914 6838 19000 6848
rect 3918 4568 4074 4668
rect 7342 4568 7498 4668
rect 10766 4568 10922 4668
rect 14190 4568 14346 4668
rect 17614 4568 17770 4668
rect 19848 4526 20018 4602
rect 19860 4510 20018 4526
rect 19860 4458 19874 4510
rect 19926 4458 20018 4510
rect 19860 4445 20018 4458
rect 19942 4432 20018 4445
rect 1754 2332 1910 2432
rect 5178 2332 5334 2432
rect 8602 2332 8758 2432
rect 12026 2332 12182 2432
rect 15450 2332 15606 2432
rect 18874 2332 19030 2432
rect 7452 146 7528 152
rect 7452 82 7458 146
rect 7522 82 7528 146
rect 7452 76 7528 82
rect 7594 146 7670 152
rect 7594 82 7600 146
rect 7664 82 7670 146
rect 7594 76 7670 82
rect 7738 146 7814 152
rect 7738 82 7744 146
rect 7808 82 7814 146
rect 7738 76 7814 82
rect 13046 146 13122 152
rect 13046 82 13052 146
rect 13116 82 13122 146
rect 13046 76 13122 82
rect 13206 146 13282 152
rect 13206 82 13212 146
rect 13276 82 13282 146
rect 13206 76 13282 82
rect 13350 146 13426 152
rect 13350 82 13356 146
rect 13420 82 13426 146
rect 13350 76 13426 82
rect 18586 146 18662 152
rect 18586 82 18592 146
rect 18656 82 18662 146
rect 18586 76 18662 82
rect 18730 146 18806 152
rect 18730 82 18736 146
rect 18800 82 18806 146
rect 18730 76 18806 82
rect 18874 146 18950 152
rect 18874 82 18880 146
rect 18944 82 18950 146
rect 18874 76 18950 82
rect 4598 -92 5062 -80
rect 4598 -168 4612 -92
rect 4688 -168 4732 -92
rect 4808 -168 4852 -92
rect 4928 -168 4972 -92
rect 5048 -168 5062 -92
rect 4598 -180 5062 -168
rect 10118 -92 10582 -80
rect 10118 -168 10132 -92
rect 10208 -168 10252 -92
rect 10328 -168 10372 -92
rect 10448 -168 10492 -92
rect 10568 -168 10582 -92
rect 10118 -180 10582 -168
rect 15758 -92 16222 -80
rect 15758 -168 15772 -92
rect 15848 -168 15892 -92
rect 15968 -168 16012 -92
rect 16088 -168 16132 -92
rect 16208 -168 16222 -92
rect 15758 -180 16222 -168
<< via1 >>
rect 4632 7164 4708 7168
rect 4632 7096 4636 7164
rect 4636 7096 4704 7164
rect 4704 7096 4708 7164
rect 4632 7092 4708 7096
rect 4752 7164 4828 7168
rect 4752 7096 4756 7164
rect 4756 7096 4824 7164
rect 4824 7096 4828 7164
rect 4752 7092 4828 7096
rect 4872 7164 4948 7168
rect 4872 7096 4876 7164
rect 4876 7096 4944 7164
rect 4944 7096 4948 7164
rect 4872 7092 4948 7096
rect 4992 7164 5068 7168
rect 4992 7096 4996 7164
rect 4996 7096 5064 7164
rect 5064 7096 5068 7164
rect 4992 7092 5068 7096
rect 10152 7164 10228 7168
rect 10152 7096 10156 7164
rect 10156 7096 10224 7164
rect 10224 7096 10228 7164
rect 10152 7092 10228 7096
rect 10272 7164 10348 7168
rect 10272 7096 10276 7164
rect 10276 7096 10344 7164
rect 10344 7096 10348 7164
rect 10272 7092 10348 7096
rect 10392 7164 10468 7168
rect 10392 7096 10396 7164
rect 10396 7096 10464 7164
rect 10464 7096 10468 7164
rect 10392 7092 10468 7096
rect 10512 7164 10588 7168
rect 10512 7096 10516 7164
rect 10516 7096 10584 7164
rect 10584 7096 10588 7164
rect 10512 7092 10588 7096
rect 15792 7164 15868 7168
rect 15792 7096 15796 7164
rect 15796 7096 15864 7164
rect 15864 7096 15868 7164
rect 15792 7092 15868 7096
rect 15912 7164 15988 7168
rect 15912 7096 15916 7164
rect 15916 7096 15984 7164
rect 15984 7096 15988 7164
rect 15912 7092 15988 7096
rect 16032 7164 16108 7168
rect 16032 7096 16036 7164
rect 16036 7096 16104 7164
rect 16104 7096 16108 7164
rect 16032 7092 16108 7096
rect 16152 7164 16228 7168
rect 16152 7096 16156 7164
rect 16156 7096 16224 7164
rect 16224 7096 16228 7164
rect 16152 7092 16228 7096
rect 1818 6854 1882 6918
rect 1960 6854 2024 6918
rect 2104 6854 2168 6918
rect 7428 6854 7492 6918
rect 7572 6854 7636 6918
rect 7716 6854 7780 6918
rect 12952 6854 13016 6918
rect 13096 6854 13160 6918
rect 13256 6854 13320 6918
rect 18564 6854 18628 6918
rect 18708 6854 18772 6918
rect 18848 6854 18912 6918
rect 19874 4504 19926 4510
rect 19874 4464 19880 4504
rect 19880 4464 19920 4504
rect 19920 4464 19926 4504
rect 19874 4458 19926 4464
rect 1760 82 1824 146
rect 1916 82 1980 146
rect 2060 82 2124 146
rect 7458 82 7522 146
rect 7600 82 7664 146
rect 7744 82 7808 146
rect 13052 82 13116 146
rect 13212 82 13276 146
rect 13356 82 13420 146
rect 18592 82 18656 146
rect 18736 82 18800 146
rect 18880 82 18944 146
rect 4612 -96 4688 -92
rect 4612 -164 4616 -96
rect 4616 -164 4684 -96
rect 4684 -164 4688 -96
rect 4612 -168 4688 -164
rect 4732 -96 4808 -92
rect 4732 -164 4736 -96
rect 4736 -164 4804 -96
rect 4804 -164 4808 -96
rect 4732 -168 4808 -164
rect 4852 -96 4928 -92
rect 4852 -164 4856 -96
rect 4856 -164 4924 -96
rect 4924 -164 4928 -96
rect 4852 -168 4928 -164
rect 4972 -96 5048 -92
rect 4972 -164 4976 -96
rect 4976 -164 5044 -96
rect 5044 -164 5048 -96
rect 4972 -168 5048 -164
rect 10132 -96 10208 -92
rect 10132 -164 10136 -96
rect 10136 -164 10204 -96
rect 10204 -164 10208 -96
rect 10132 -168 10208 -164
rect 10252 -96 10328 -92
rect 10252 -164 10256 -96
rect 10256 -164 10324 -96
rect 10324 -164 10328 -96
rect 10252 -168 10328 -164
rect 10372 -96 10448 -92
rect 10372 -164 10376 -96
rect 10376 -164 10444 -96
rect 10444 -164 10448 -96
rect 10372 -168 10448 -164
rect 10492 -96 10568 -92
rect 10492 -164 10496 -96
rect 10496 -164 10564 -96
rect 10564 -164 10568 -96
rect 10492 -168 10568 -164
rect 15772 -96 15848 -92
rect 15772 -164 15776 -96
rect 15776 -164 15844 -96
rect 15844 -164 15848 -96
rect 15772 -168 15848 -164
rect 15892 -96 15968 -92
rect 15892 -164 15896 -96
rect 15896 -164 15964 -96
rect 15964 -164 15968 -96
rect 15892 -168 15968 -164
rect 16012 -96 16088 -92
rect 16012 -164 16016 -96
rect 16016 -164 16084 -96
rect 16084 -164 16088 -96
rect 16012 -168 16088 -164
rect 16132 -96 16208 -92
rect 16132 -164 16136 -96
rect 16136 -164 16204 -96
rect 16204 -164 16208 -96
rect 16132 -168 16208 -164
<< metal2 >>
rect 4618 7172 5082 7180
rect 4618 7088 4628 7172
rect 4712 7088 4748 7172
rect 4832 7088 4868 7172
rect 4952 7088 4988 7172
rect 5072 7088 5082 7172
rect 4618 7080 5082 7088
rect 10138 7172 10602 7180
rect 10138 7088 10148 7172
rect 10232 7088 10268 7172
rect 10352 7088 10388 7172
rect 10472 7088 10508 7172
rect 10592 7088 10602 7172
rect 10138 7080 10602 7088
rect 15778 7172 16242 7180
rect 15778 7088 15788 7172
rect 15872 7088 15908 7172
rect 15992 7088 16028 7172
rect 16112 7088 16148 7172
rect 16232 7088 16242 7172
rect 15778 7080 16242 7088
rect 1804 6922 1896 6932
rect 1804 6850 1814 6922
rect 1886 6850 1896 6922
rect 1804 6840 1896 6850
rect 1946 6922 2038 6932
rect 1946 6850 1956 6922
rect 2028 6850 2038 6922
rect 1946 6840 2038 6850
rect 2090 6922 2182 6932
rect 2090 6850 2100 6922
rect 2172 6850 2182 6922
rect 2090 6840 2182 6850
rect 7414 6922 7506 6932
rect 7414 6850 7424 6922
rect 7496 6850 7506 6922
rect 7414 6840 7506 6850
rect 7558 6922 7650 6932
rect 7558 6850 7568 6922
rect 7640 6850 7650 6922
rect 7558 6840 7650 6850
rect 7702 6922 7794 6932
rect 7702 6850 7712 6922
rect 7784 6850 7794 6922
rect 7702 6840 7794 6850
rect 12938 6922 13030 6932
rect 12938 6850 12948 6922
rect 13020 6850 13030 6922
rect 12938 6840 13030 6850
rect 13082 6922 13174 6932
rect 13082 6850 13092 6922
rect 13164 6850 13174 6922
rect 13082 6840 13174 6850
rect 13242 6922 13334 6932
rect 13242 6850 13252 6922
rect 13324 6850 13334 6922
rect 13242 6840 13334 6850
rect 18550 6922 18642 6932
rect 18550 6850 18560 6922
rect 18632 6850 18642 6922
rect 18550 6840 18642 6850
rect 18694 6922 18786 6932
rect 18694 6850 18704 6922
rect 18776 6850 18786 6922
rect 18694 6840 18786 6850
rect 18834 6922 18926 6932
rect 18834 6850 18844 6922
rect 18916 6850 18926 6922
rect 18834 6840 18926 6850
rect 19848 4526 20018 4602
rect 19860 4512 20018 4526
rect 19860 4456 19872 4512
rect 19928 4456 20018 4512
rect 19860 4445 20018 4456
rect 19942 4432 20018 4445
rect 1746 150 1838 160
rect 1746 78 1756 150
rect 1828 78 1838 150
rect 1746 68 1838 78
rect 1902 150 1994 160
rect 1902 78 1912 150
rect 1984 78 1994 150
rect 1902 68 1994 78
rect 2046 150 2138 160
rect 2046 78 2056 150
rect 2128 78 2138 150
rect 2046 68 2138 78
rect 7444 150 7536 160
rect 7444 78 7454 150
rect 7526 78 7536 150
rect 7444 68 7536 78
rect 7586 150 7678 160
rect 7586 78 7596 150
rect 7668 78 7678 150
rect 7586 68 7678 78
rect 7730 150 7822 160
rect 7730 78 7740 150
rect 7812 78 7822 150
rect 7730 68 7822 78
rect 13038 150 13130 160
rect 13038 78 13048 150
rect 13120 78 13130 150
rect 13038 68 13130 78
rect 13198 150 13290 160
rect 13198 78 13208 150
rect 13280 78 13290 150
rect 13198 68 13290 78
rect 13342 150 13434 160
rect 13342 78 13352 150
rect 13424 78 13434 150
rect 13342 68 13434 78
rect 18578 150 18670 160
rect 18578 78 18588 150
rect 18660 78 18670 150
rect 18578 68 18670 78
rect 18722 150 18814 160
rect 18722 78 18732 150
rect 18804 78 18814 150
rect 18722 68 18814 78
rect 18866 150 18958 160
rect 18866 78 18876 150
rect 18948 78 18958 150
rect 18866 68 18958 78
rect 4598 -88 5062 -80
rect 4598 -172 4608 -88
rect 4692 -172 4728 -88
rect 4812 -172 4848 -88
rect 4932 -172 4968 -88
rect 5052 -172 5062 -88
rect 4598 -180 5062 -172
rect 10118 -88 10582 -80
rect 10118 -172 10128 -88
rect 10212 -172 10248 -88
rect 10332 -172 10368 -88
rect 10452 -172 10488 -88
rect 10572 -172 10582 -88
rect 10118 -180 10582 -172
rect 15758 -88 16222 -80
rect 15758 -172 15768 -88
rect 15852 -172 15888 -88
rect 15972 -172 16008 -88
rect 16092 -172 16128 -88
rect 16212 -172 16222 -88
rect 15758 -180 16222 -172
<< via2 >>
rect 4628 7168 4712 7172
rect 4628 7092 4632 7168
rect 4632 7092 4708 7168
rect 4708 7092 4712 7168
rect 4628 7088 4712 7092
rect 4748 7168 4832 7172
rect 4748 7092 4752 7168
rect 4752 7092 4828 7168
rect 4828 7092 4832 7168
rect 4748 7088 4832 7092
rect 4868 7168 4952 7172
rect 4868 7092 4872 7168
rect 4872 7092 4948 7168
rect 4948 7092 4952 7168
rect 4868 7088 4952 7092
rect 4988 7168 5072 7172
rect 4988 7092 4992 7168
rect 4992 7092 5068 7168
rect 5068 7092 5072 7168
rect 4988 7088 5072 7092
rect 10148 7168 10232 7172
rect 10148 7092 10152 7168
rect 10152 7092 10228 7168
rect 10228 7092 10232 7168
rect 10148 7088 10232 7092
rect 10268 7168 10352 7172
rect 10268 7092 10272 7168
rect 10272 7092 10348 7168
rect 10348 7092 10352 7168
rect 10268 7088 10352 7092
rect 10388 7168 10472 7172
rect 10388 7092 10392 7168
rect 10392 7092 10468 7168
rect 10468 7092 10472 7168
rect 10388 7088 10472 7092
rect 10508 7168 10592 7172
rect 10508 7092 10512 7168
rect 10512 7092 10588 7168
rect 10588 7092 10592 7168
rect 10508 7088 10592 7092
rect 15788 7168 15872 7172
rect 15788 7092 15792 7168
rect 15792 7092 15868 7168
rect 15868 7092 15872 7168
rect 15788 7088 15872 7092
rect 15908 7168 15992 7172
rect 15908 7092 15912 7168
rect 15912 7092 15988 7168
rect 15988 7092 15992 7168
rect 15908 7088 15992 7092
rect 16028 7168 16112 7172
rect 16028 7092 16032 7168
rect 16032 7092 16108 7168
rect 16108 7092 16112 7168
rect 16028 7088 16112 7092
rect 16148 7168 16232 7172
rect 16148 7092 16152 7168
rect 16152 7092 16228 7168
rect 16228 7092 16232 7168
rect 16148 7088 16232 7092
rect 1814 6918 1886 6922
rect 1814 6854 1818 6918
rect 1818 6854 1882 6918
rect 1882 6854 1886 6918
rect 1814 6850 1886 6854
rect 1956 6918 2028 6922
rect 1956 6854 1960 6918
rect 1960 6854 2024 6918
rect 2024 6854 2028 6918
rect 1956 6850 2028 6854
rect 2100 6918 2172 6922
rect 2100 6854 2104 6918
rect 2104 6854 2168 6918
rect 2168 6854 2172 6918
rect 2100 6850 2172 6854
rect 7424 6918 7496 6922
rect 7424 6854 7428 6918
rect 7428 6854 7492 6918
rect 7492 6854 7496 6918
rect 7424 6850 7496 6854
rect 7568 6918 7640 6922
rect 7568 6854 7572 6918
rect 7572 6854 7636 6918
rect 7636 6854 7640 6918
rect 7568 6850 7640 6854
rect 7712 6918 7784 6922
rect 7712 6854 7716 6918
rect 7716 6854 7780 6918
rect 7780 6854 7784 6918
rect 7712 6850 7784 6854
rect 12948 6918 13020 6922
rect 12948 6854 12952 6918
rect 12952 6854 13016 6918
rect 13016 6854 13020 6918
rect 12948 6850 13020 6854
rect 13092 6918 13164 6922
rect 13092 6854 13096 6918
rect 13096 6854 13160 6918
rect 13160 6854 13164 6918
rect 13092 6850 13164 6854
rect 13252 6918 13324 6922
rect 13252 6854 13256 6918
rect 13256 6854 13320 6918
rect 13320 6854 13324 6918
rect 13252 6850 13324 6854
rect 18560 6918 18632 6922
rect 18560 6854 18564 6918
rect 18564 6854 18628 6918
rect 18628 6854 18632 6918
rect 18560 6850 18632 6854
rect 18704 6918 18776 6922
rect 18704 6854 18708 6918
rect 18708 6854 18772 6918
rect 18772 6854 18776 6918
rect 18704 6850 18776 6854
rect 18844 6918 18916 6922
rect 18844 6854 18848 6918
rect 18848 6854 18912 6918
rect 18912 6854 18916 6918
rect 18844 6850 18916 6854
rect 19872 4510 19928 4512
rect 19872 4458 19874 4510
rect 19874 4458 19926 4510
rect 19926 4458 19928 4510
rect 19872 4456 19928 4458
rect 1756 146 1828 150
rect 1756 82 1760 146
rect 1760 82 1824 146
rect 1824 82 1828 146
rect 1756 78 1828 82
rect 1912 146 1984 150
rect 1912 82 1916 146
rect 1916 82 1980 146
rect 1980 82 1984 146
rect 1912 78 1984 82
rect 2056 146 2128 150
rect 2056 82 2060 146
rect 2060 82 2124 146
rect 2124 82 2128 146
rect 2056 78 2128 82
rect 7454 146 7526 150
rect 7454 82 7458 146
rect 7458 82 7522 146
rect 7522 82 7526 146
rect 7454 78 7526 82
rect 7596 146 7668 150
rect 7596 82 7600 146
rect 7600 82 7664 146
rect 7664 82 7668 146
rect 7596 78 7668 82
rect 7740 146 7812 150
rect 7740 82 7744 146
rect 7744 82 7808 146
rect 7808 82 7812 146
rect 7740 78 7812 82
rect 13048 146 13120 150
rect 13048 82 13052 146
rect 13052 82 13116 146
rect 13116 82 13120 146
rect 13048 78 13120 82
rect 13208 146 13280 150
rect 13208 82 13212 146
rect 13212 82 13276 146
rect 13276 82 13280 146
rect 13208 78 13280 82
rect 13352 146 13424 150
rect 13352 82 13356 146
rect 13356 82 13420 146
rect 13420 82 13424 146
rect 13352 78 13424 82
rect 18588 146 18660 150
rect 18588 82 18592 146
rect 18592 82 18656 146
rect 18656 82 18660 146
rect 18588 78 18660 82
rect 18732 146 18804 150
rect 18732 82 18736 146
rect 18736 82 18800 146
rect 18800 82 18804 146
rect 18732 78 18804 82
rect 18876 146 18948 150
rect 18876 82 18880 146
rect 18880 82 18944 146
rect 18944 82 18948 146
rect 18876 78 18948 82
rect 4608 -92 4692 -88
rect 4608 -168 4612 -92
rect 4612 -168 4688 -92
rect 4688 -168 4692 -92
rect 4608 -172 4692 -168
rect 4728 -92 4812 -88
rect 4728 -168 4732 -92
rect 4732 -168 4808 -92
rect 4808 -168 4812 -92
rect 4728 -172 4812 -168
rect 4848 -92 4932 -88
rect 4848 -168 4852 -92
rect 4852 -168 4928 -92
rect 4928 -168 4932 -92
rect 4848 -172 4932 -168
rect 4968 -92 5052 -88
rect 4968 -168 4972 -92
rect 4972 -168 5048 -92
rect 5048 -168 5052 -92
rect 4968 -172 5052 -168
rect 10128 -92 10212 -88
rect 10128 -168 10132 -92
rect 10132 -168 10208 -92
rect 10208 -168 10212 -92
rect 10128 -172 10212 -168
rect 10248 -92 10332 -88
rect 10248 -168 10252 -92
rect 10252 -168 10328 -92
rect 10328 -168 10332 -92
rect 10248 -172 10332 -168
rect 10368 -92 10452 -88
rect 10368 -168 10372 -92
rect 10372 -168 10448 -92
rect 10448 -168 10452 -92
rect 10368 -172 10452 -168
rect 10488 -92 10572 -88
rect 10488 -168 10492 -92
rect 10492 -168 10568 -92
rect 10568 -168 10572 -92
rect 10488 -172 10572 -168
rect 15768 -92 15852 -88
rect 15768 -168 15772 -92
rect 15772 -168 15848 -92
rect 15848 -168 15852 -92
rect 15768 -172 15852 -168
rect 15888 -92 15972 -88
rect 15888 -168 15892 -92
rect 15892 -168 15968 -92
rect 15968 -168 15972 -92
rect 15888 -172 15972 -168
rect 16008 -92 16092 -88
rect 16008 -168 16012 -92
rect 16012 -168 16088 -92
rect 16088 -168 16092 -92
rect 16008 -172 16092 -168
rect 16128 -92 16212 -88
rect 16128 -168 16132 -92
rect 16132 -168 16208 -92
rect 16208 -168 16212 -92
rect 16128 -172 16212 -168
<< metal3 >>
rect 4618 7176 5082 7180
rect 4618 7084 4624 7176
rect 4716 7084 4744 7176
rect 4836 7084 4864 7176
rect 4956 7084 4984 7176
rect 5076 7084 5082 7176
rect 4618 7080 5082 7084
rect 10138 7176 10602 7180
rect 10138 7084 10144 7176
rect 10236 7084 10264 7176
rect 10356 7084 10384 7176
rect 10476 7084 10504 7176
rect 10596 7084 10602 7176
rect 10138 7080 10602 7084
rect 15778 7176 16242 7180
rect 15778 7084 15784 7176
rect 15876 7084 15904 7176
rect 15996 7084 16024 7176
rect 16116 7084 16144 7176
rect 16236 7084 16242 7176
rect 15778 7080 16242 7084
rect 1800 6932 2170 6938
rect 1800 6926 2182 6932
rect 1800 6846 1810 6926
rect 1890 6846 1952 6926
rect 2032 6846 2096 6926
rect 2176 6846 2182 6926
rect 1800 6840 2182 6846
rect 7412 6926 7796 6938
rect 7412 6846 7420 6926
rect 7500 6846 7564 6926
rect 7644 6846 7708 6926
rect 7788 6846 7796 6926
rect 1800 6838 2170 6840
rect 7412 6838 7796 6846
rect 12936 6926 13336 6938
rect 12936 6846 12944 6926
rect 13024 6846 13088 6926
rect 13168 6846 13248 6926
rect 13328 6846 13336 6926
rect 12936 6838 13336 6846
rect 18548 6926 18932 6938
rect 18548 6846 18556 6926
rect 18636 6846 18700 6926
rect 18780 6846 18840 6926
rect 18920 6846 18932 6926
rect 18548 6838 18932 6846
rect 19702 4512 20018 4602
rect 19702 4456 19872 4512
rect 19928 4456 20018 4512
rect 19702 3601 20018 4456
rect 1746 154 2138 162
rect 1746 74 1752 154
rect 1832 74 1908 154
rect 1988 74 2052 154
rect 2132 74 2138 154
rect 1746 62 2138 74
rect 7442 154 7826 162
rect 7442 74 7450 154
rect 7530 74 7592 154
rect 7672 74 7736 154
rect 7816 74 7826 154
rect 7442 62 7826 74
rect 13036 154 13436 162
rect 13036 74 13044 154
rect 13124 74 13204 154
rect 13284 74 13348 154
rect 13428 74 13436 154
rect 13036 62 13436 74
rect 18576 154 18960 162
rect 18576 74 18584 154
rect 18664 74 18728 154
rect 18808 74 18872 154
rect 18952 74 18960 154
rect 18576 62 18960 74
rect 4598 -84 5062 -80
rect 4598 -176 4604 -84
rect 4696 -176 4724 -84
rect 4816 -176 4844 -84
rect 4936 -176 4964 -84
rect 5056 -176 5062 -84
rect 4598 -180 5062 -176
rect 10118 -84 10582 -80
rect 10118 -176 10124 -84
rect 10216 -176 10244 -84
rect 10336 -176 10364 -84
rect 10456 -176 10484 -84
rect 10576 -176 10582 -84
rect 10118 -180 10582 -176
rect 15758 -84 16222 -80
rect 15758 -176 15764 -84
rect 15856 -176 15884 -84
rect 15976 -176 16004 -84
rect 16096 -176 16124 -84
rect 16216 -176 16222 -84
rect 15758 -180 16222 -176
<< via3 >>
rect 4624 7172 4716 7176
rect 4624 7088 4628 7172
rect 4628 7088 4712 7172
rect 4712 7088 4716 7172
rect 4624 7084 4716 7088
rect 4744 7172 4836 7176
rect 4744 7088 4748 7172
rect 4748 7088 4832 7172
rect 4832 7088 4836 7172
rect 4744 7084 4836 7088
rect 4864 7172 4956 7176
rect 4864 7088 4868 7172
rect 4868 7088 4952 7172
rect 4952 7088 4956 7172
rect 4864 7084 4956 7088
rect 4984 7172 5076 7176
rect 4984 7088 4988 7172
rect 4988 7088 5072 7172
rect 5072 7088 5076 7172
rect 4984 7084 5076 7088
rect 10144 7172 10236 7176
rect 10144 7088 10148 7172
rect 10148 7088 10232 7172
rect 10232 7088 10236 7172
rect 10144 7084 10236 7088
rect 10264 7172 10356 7176
rect 10264 7088 10268 7172
rect 10268 7088 10352 7172
rect 10352 7088 10356 7172
rect 10264 7084 10356 7088
rect 10384 7172 10476 7176
rect 10384 7088 10388 7172
rect 10388 7088 10472 7172
rect 10472 7088 10476 7172
rect 10384 7084 10476 7088
rect 10504 7172 10596 7176
rect 10504 7088 10508 7172
rect 10508 7088 10592 7172
rect 10592 7088 10596 7172
rect 10504 7084 10596 7088
rect 15784 7172 15876 7176
rect 15784 7088 15788 7172
rect 15788 7088 15872 7172
rect 15872 7088 15876 7172
rect 15784 7084 15876 7088
rect 15904 7172 15996 7176
rect 15904 7088 15908 7172
rect 15908 7088 15992 7172
rect 15992 7088 15996 7172
rect 15904 7084 15996 7088
rect 16024 7172 16116 7176
rect 16024 7088 16028 7172
rect 16028 7088 16112 7172
rect 16112 7088 16116 7172
rect 16024 7084 16116 7088
rect 16144 7172 16236 7176
rect 16144 7088 16148 7172
rect 16148 7088 16232 7172
rect 16232 7088 16236 7172
rect 16144 7084 16236 7088
rect 1810 6922 1890 6926
rect 1810 6850 1814 6922
rect 1814 6850 1886 6922
rect 1886 6850 1890 6922
rect 1810 6846 1890 6850
rect 1952 6922 2032 6926
rect 1952 6850 1956 6922
rect 1956 6850 2028 6922
rect 2028 6850 2032 6922
rect 1952 6846 2032 6850
rect 2096 6922 2176 6926
rect 2096 6850 2100 6922
rect 2100 6850 2172 6922
rect 2172 6850 2176 6922
rect 2096 6846 2176 6850
rect 7420 6922 7500 6926
rect 7420 6850 7424 6922
rect 7424 6850 7496 6922
rect 7496 6850 7500 6922
rect 7420 6846 7500 6850
rect 7564 6922 7644 6926
rect 7564 6850 7568 6922
rect 7568 6850 7640 6922
rect 7640 6850 7644 6922
rect 7564 6846 7644 6850
rect 7708 6922 7788 6926
rect 7708 6850 7712 6922
rect 7712 6850 7784 6922
rect 7784 6850 7788 6922
rect 7708 6846 7788 6850
rect 12944 6922 13024 6926
rect 12944 6850 12948 6922
rect 12948 6850 13020 6922
rect 13020 6850 13024 6922
rect 12944 6846 13024 6850
rect 13088 6922 13168 6926
rect 13088 6850 13092 6922
rect 13092 6850 13164 6922
rect 13164 6850 13168 6922
rect 13088 6846 13168 6850
rect 13248 6922 13328 6926
rect 13248 6850 13252 6922
rect 13252 6850 13324 6922
rect 13324 6850 13328 6922
rect 13248 6846 13328 6850
rect 18556 6922 18636 6926
rect 18556 6850 18560 6922
rect 18560 6850 18632 6922
rect 18632 6850 18636 6922
rect 18556 6846 18636 6850
rect 18700 6922 18780 6926
rect 18700 6850 18704 6922
rect 18704 6850 18776 6922
rect 18776 6850 18780 6922
rect 18700 6846 18780 6850
rect 18840 6922 18920 6926
rect 18840 6850 18844 6922
rect 18844 6850 18916 6922
rect 18916 6850 18920 6922
rect 18840 6846 18920 6850
rect 1752 150 1832 154
rect 1752 78 1756 150
rect 1756 78 1828 150
rect 1828 78 1832 150
rect 1752 74 1832 78
rect 1908 150 1988 154
rect 1908 78 1912 150
rect 1912 78 1984 150
rect 1984 78 1988 150
rect 1908 74 1988 78
rect 2052 150 2132 154
rect 2052 78 2056 150
rect 2056 78 2128 150
rect 2128 78 2132 150
rect 2052 74 2132 78
rect 7450 150 7530 154
rect 7450 78 7454 150
rect 7454 78 7526 150
rect 7526 78 7530 150
rect 7450 74 7530 78
rect 7592 150 7672 154
rect 7592 78 7596 150
rect 7596 78 7668 150
rect 7668 78 7672 150
rect 7592 74 7672 78
rect 7736 150 7816 154
rect 7736 78 7740 150
rect 7740 78 7812 150
rect 7812 78 7816 150
rect 7736 74 7816 78
rect 13044 150 13124 154
rect 13044 78 13048 150
rect 13048 78 13120 150
rect 13120 78 13124 150
rect 13044 74 13124 78
rect 13204 150 13284 154
rect 13204 78 13208 150
rect 13208 78 13280 150
rect 13280 78 13284 150
rect 13204 74 13284 78
rect 13348 150 13428 154
rect 13348 78 13352 150
rect 13352 78 13424 150
rect 13424 78 13428 150
rect 13348 74 13428 78
rect 18584 150 18664 154
rect 18584 78 18588 150
rect 18588 78 18660 150
rect 18660 78 18664 150
rect 18584 74 18664 78
rect 18728 150 18808 154
rect 18728 78 18732 150
rect 18732 78 18804 150
rect 18804 78 18808 150
rect 18728 74 18808 78
rect 18872 150 18952 154
rect 18872 78 18876 150
rect 18876 78 18948 150
rect 18948 78 18952 150
rect 18872 74 18952 78
rect 4604 -88 4696 -84
rect 4604 -172 4608 -88
rect 4608 -172 4692 -88
rect 4692 -172 4696 -88
rect 4604 -176 4696 -172
rect 4724 -88 4816 -84
rect 4724 -172 4728 -88
rect 4728 -172 4812 -88
rect 4812 -172 4816 -88
rect 4724 -176 4816 -172
rect 4844 -88 4936 -84
rect 4844 -172 4848 -88
rect 4848 -172 4932 -88
rect 4932 -172 4936 -88
rect 4844 -176 4936 -172
rect 4964 -88 5056 -84
rect 4964 -172 4968 -88
rect 4968 -172 5052 -88
rect 5052 -172 5056 -88
rect 4964 -176 5056 -172
rect 10124 -88 10216 -84
rect 10124 -172 10128 -88
rect 10128 -172 10212 -88
rect 10212 -172 10216 -88
rect 10124 -176 10216 -172
rect 10244 -88 10336 -84
rect 10244 -172 10248 -88
rect 10248 -172 10332 -88
rect 10332 -172 10336 -88
rect 10244 -176 10336 -172
rect 10364 -88 10456 -84
rect 10364 -172 10368 -88
rect 10368 -172 10452 -88
rect 10452 -172 10456 -88
rect 10364 -176 10456 -172
rect 10484 -88 10576 -84
rect 10484 -172 10488 -88
rect 10488 -172 10572 -88
rect 10572 -172 10576 -88
rect 10484 -176 10576 -172
rect 15764 -88 15856 -84
rect 15764 -172 15768 -88
rect 15768 -172 15852 -88
rect 15852 -172 15856 -88
rect 15764 -176 15856 -172
rect 15884 -88 15976 -84
rect 15884 -172 15888 -88
rect 15888 -172 15972 -88
rect 15972 -172 15976 -88
rect 15884 -176 15976 -172
rect 16004 -88 16096 -84
rect 16004 -172 16008 -88
rect 16008 -172 16092 -88
rect 16092 -172 16096 -88
rect 16004 -176 16096 -172
rect 16124 -88 16216 -84
rect 16124 -172 16128 -88
rect 16128 -172 16212 -88
rect 16212 -172 16216 -88
rect 16124 -176 16216 -172
<< metal4 >>
rect 4618 7176 5082 7180
rect 4618 7084 4624 7176
rect 4716 7084 4744 7176
rect 4836 7084 4864 7176
rect 4956 7084 4984 7176
rect 5076 7084 5082 7176
rect 4618 7080 5082 7084
rect 10138 7176 10250 7180
rect 10138 7084 10144 7176
rect 10236 7084 10250 7176
rect 10138 7080 10250 7084
rect 10600 7080 10602 7180
rect 15778 7176 16242 7180
rect 15778 7084 15784 7176
rect 15876 7084 15904 7176
rect 15996 7084 16024 7176
rect 16116 7084 16144 7176
rect 16236 7084 16242 7176
rect 15778 7080 16242 7084
rect 7412 6926 7508 6938
rect 7412 6846 7420 6926
rect 7500 6846 7508 6926
rect 7412 6838 7508 6846
rect 7556 6926 7652 6938
rect 7556 6846 7564 6926
rect 7644 6846 7652 6926
rect 7556 6838 7652 6846
rect 7700 6926 7796 6938
rect 7700 6846 7708 6926
rect 7788 6846 7796 6926
rect 7700 6838 7796 6846
rect 12936 6926 13032 6938
rect 12936 6846 12944 6926
rect 13024 6846 13032 6926
rect 12936 6838 13032 6846
rect 13080 6926 13176 6938
rect 13080 6846 13088 6926
rect 13168 6846 13176 6926
rect 13080 6838 13176 6846
rect 13240 6926 13336 6938
rect 13240 6846 13248 6926
rect 13328 6846 13336 6926
rect 13240 6838 13336 6846
rect 18548 6926 18644 6938
rect 18548 6846 18556 6926
rect 18636 6846 18644 6926
rect 18548 6838 18644 6846
rect 18692 6926 18788 6938
rect 18692 6846 18700 6926
rect 18780 6846 18788 6926
rect 18692 6838 18788 6846
rect 18832 6926 18928 6938
rect 18832 6846 18840 6926
rect 18920 6846 18928 6926
rect 18832 6838 18928 6846
rect 1746 154 2138 162
rect 1746 74 1752 154
rect 1832 74 1908 154
rect 1988 74 2052 154
rect 2132 74 2138 154
rect 1746 62 2138 74
rect 7442 154 7538 162
rect 7442 74 7450 154
rect 7530 74 7538 154
rect 7442 62 7538 74
rect 7584 154 7680 162
rect 7584 74 7592 154
rect 7672 74 7680 154
rect 7584 62 7680 74
rect 7728 154 7824 162
rect 7728 74 7736 154
rect 7816 74 7824 154
rect 7728 62 7824 74
rect 13036 154 13132 162
rect 13036 74 13044 154
rect 13124 74 13132 154
rect 13036 62 13132 74
rect 13196 154 13292 162
rect 13196 74 13204 154
rect 13284 74 13292 154
rect 13196 62 13292 74
rect 13340 154 13436 162
rect 13340 74 13348 154
rect 13428 74 13436 154
rect 13340 62 13436 74
rect 18576 154 18672 162
rect 18576 74 18584 154
rect 18664 74 18672 154
rect 18576 62 18672 74
rect 18720 154 18816 162
rect 18720 74 18728 154
rect 18808 74 18816 154
rect 18720 62 18816 74
rect 18864 154 18960 162
rect 18864 74 18872 154
rect 18952 74 18960 154
rect 18864 62 18960 74
rect 4598 -84 5062 -80
rect 4598 -176 4604 -84
rect 4696 -176 4724 -84
rect 4816 -176 4844 -84
rect 4936 -176 4964 -84
rect 5056 -176 5062 -84
rect 4598 -180 5062 -176
rect 10118 -84 10582 -80
rect 10118 -176 10124 -84
rect 10216 -176 10244 -84
rect 10336 -176 10364 -84
rect 10456 -176 10484 -84
rect 10576 -176 10582 -84
rect 10118 -180 10582 -176
rect 15758 -84 16222 -80
rect 15758 -176 15764 -84
rect 15856 -176 15884 -84
rect 15976 -176 16004 -84
rect 16096 -176 16124 -84
rect 16216 -176 16222 -84
rect 15758 -180 16222 -176
use res_pdiff  res_pdiff_1
timestamp 1637571367
transform 0 1 19836 -1 0 4684
box 0 0 450 900
use res_pdiff  res_pdiff_0
timestamp 1637571367
transform 1 0 19620 0 1 4420
box 0 0 450 900
use ring_osc  ring_osc_0
timestamp 1637401559
transform 1 0 600 0 1 62
box -600 -62 21100 6938
use pwell_co_ring  pwell_co_ring_0
timestamp 1637401559
transform 1 0 340 0 1 -160
box 0 0 21120 7320
use power_ring  power_ring_0
timestamp 1637401559
transform 1 0 -1800 0 1 -7000
box 0 0 24400 21000
<< labels >>
flabel metal1 1824 2382 1824 2382 1 FreeSans 1600 0 0 0 p[0]
port 1 s signal output
flabel metal1 5248 2382 5248 2382 1 FreeSans 1600 0 0 0 p[2]
port 3 s signal output
flabel metal1 8672 2382 8672 2382 1 FreeSans 1600 0 0 0 p[4]
port 5 s signal output
flabel metal1 12096 2382 12096 2382 1 FreeSans 1600 0 0 0 p[6]
port 7 s signal output
flabel metal1 15520 2382 15520 2382 1 FreeSans 1600 0 0 0 p[8]
port 9 s signal output
flabel metal1 18944 2382 18944 2382 1 FreeSans 1600 0 0 0 p[10]
port 11 s signal output
flabel metal1 4004 4618 4004 4618 1 FreeSans 1600 0 0 0 p[1]
port 2 s signal output
flabel metal1 7428 4618 7428 4618 1 FreeSans 1600 0 0 0 p[3]
port 4 s signal output
flabel metal1 10852 4618 10852 4618 1 FreeSans 1600 0 0 0 p[5]
port 6 s signal output
flabel metal1 14276 4618 14276 4618 1 FreeSans 1600 0 0 0 p[7]
port 8 s signal output
flabel metal1 17700 4618 17700 4618 1 FreeSans 1600 0 0 0 p[9]
port 10 s signal output
<< end >>
