magic
tech sky130A
magscale 1 2
timestamp 1624647652
<< ndiff >>
rect 1627 12258 1661 12292
<< pdiff >>
rect 1627 12582 1661 12616
<< locali >>
rect 1910 12548 1955 12592
rect 2308 12542 2353 12586
rect 62 12438 158 12460
rect 62 12382 74 12438
rect 130 12406 158 12438
rect 130 12382 142 12406
rect 1496 12384 1521 12418
rect 62 12360 142 12382
<< viali >>
rect 74 12382 130 12438
<< metal1 >>
rect 0 12656 1994 12752
rect 62 12438 142 12484
rect 62 12382 74 12438
rect 130 12382 142 12438
rect 21722 12404 23600 12476
rect 62 12348 142 12382
rect 800 12112 1962 12208
<< metal2 >>
rect 5382 13970 5566 13986
rect 5382 13910 5444 13970
rect 5504 13910 5566 13970
rect 5382 13894 5566 13910
rect 10258 13970 10442 13986
rect 10258 13910 10320 13970
rect 10380 13910 10442 13970
rect 10258 13894 10442 13910
rect 13570 13970 13754 13986
rect 13570 13910 13632 13970
rect 13692 13910 13754 13970
rect 13570 13894 13754 13910
rect 16698 13970 16882 13986
rect 16698 13910 16760 13970
rect 16820 13910 16882 13970
rect 16698 13894 16882 13910
rect 21114 13970 21298 13986
rect 21114 13910 21176 13970
rect 21236 13910 21298 13970
rect 21114 13894 21298 13910
rect 24426 11522 24610 11542
rect 24426 11462 24488 11522
rect 24548 11462 24610 11522
rect 24426 11442 24610 11462
rect 1334 7306 1518 7322
rect 1334 7246 1396 7306
rect 1456 7246 1518 7306
rect 1334 7230 1518 7246
rect 5014 7306 5198 7322
rect 5014 7246 5076 7306
rect 5136 7246 5198 7306
rect 5014 7230 5198 7246
rect 8510 7306 8694 7322
rect 8510 7246 8572 7306
rect 8632 7246 8694 7306
rect 8510 7230 8694 7246
rect 13110 7306 13294 7322
rect 13110 7246 13172 7306
rect 13232 7246 13294 7306
rect 13110 7230 13294 7246
rect 15778 7306 15962 7322
rect 15778 7246 15840 7306
rect 15900 7246 15962 7306
rect 15778 7230 15962 7246
rect 19182 7306 19366 7322
rect 19182 7246 19244 7306
rect 19304 7246 19366 7306
rect 19182 7230 19366 7246
<< via2 >>
rect 5444 13910 5504 13970
rect 10320 13910 10380 13970
rect 13632 13910 13692 13970
rect 16760 13910 16820 13970
rect 21176 13910 21236 13970
rect 24488 11462 24548 11522
rect 1396 7246 1456 7306
rect 5076 7246 5136 7306
rect 8572 7246 8632 7306
rect 13172 7246 13232 7306
rect 15840 7246 15900 7306
rect 19244 7246 19304 7306
<< metal3 >>
rect 0 20600 5200 21000
rect 5428 13970 5520 14076
rect 5428 13910 5444 13970
rect 5504 13910 5520 13970
rect 5428 13804 5520 13910
rect 10304 13970 10396 14076
rect 10304 13910 10320 13970
rect 10380 13910 10396 13970
rect 10304 13804 10396 13910
rect 13616 13970 13708 14076
rect 13616 13910 13632 13970
rect 13692 13910 13708 13970
rect 13616 13804 13708 13910
rect 16744 13970 16836 14076
rect 16744 13910 16760 13970
rect 16820 13910 16836 13970
rect 16744 13804 16836 13910
rect 21160 13970 21252 14076
rect 21160 13910 21176 13970
rect 21236 13910 21252 13970
rect 21160 13804 21252 13910
rect 24464 11522 24572 11628
rect 24464 11462 24488 11522
rect 24548 11462 24572 11522
rect 24464 11356 24572 11462
rect 1380 7306 1472 7412
rect 1380 7246 1396 7306
rect 1456 7246 1472 7306
rect 1380 7140 1472 7246
rect 5060 7306 5152 7412
rect 5060 7246 5076 7306
rect 5136 7246 5152 7306
rect 5060 7140 5152 7246
rect 8556 7306 8648 7412
rect 8556 7246 8572 7306
rect 8632 7246 8648 7306
rect 8556 7140 8648 7246
rect 13156 7306 13248 7412
rect 13156 7246 13172 7306
rect 13232 7246 13248 7306
rect 13156 7140 13248 7246
rect 15824 7306 15916 7412
rect 15824 7246 15840 7306
rect 15900 7246 15916 7306
rect 15824 7140 15916 7246
rect 19228 7306 19320 7412
rect 19228 7246 19244 7306
rect 19304 7246 19320 7306
rect 19228 7140 19320 7246
rect 18600 800 23600 1200
use ring_osc  ring_osc_0
timestamp 1624647281
transform 1 0 1500 0 1 7600
box -1410 -344 23110 6300
use via_m1  via_m1_4
timestamp 1623561200
transform 1 0 -7298 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_5
timestamp 1623561200
transform 1 0 -1698 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_8
timestamp 1623561200
transform 1 0 3902 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_9
timestamp 1623561200
transform 1 0 9502 0 1 662
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_4
timestamp 1623563441
transform 1 0 6400 0 1 7360
box 0 2 400 98
use via_m4_li  via_m4_li_5
timestamp 1623563441
transform 1 0 12000 0 1 7360
box 0 2 400 98
use pwell_co_ring  pwell_co_ring_0
timestamp 1623529308
transform 1 0 3020 0 1 13740
box -1680 -6360 20145 60
use via_m1  via_m1_3
timestamp 1623561200
transform 1 0 -7298 0 1 6498
box 10898 6956 11298 7052
use via_m1  via_m1_2
timestamp 1623561200
transform 1 0 -10098 0 1 5156
box 10898 6956 11298 7052
use via_m1  via_m1_1
timestamp 1623561200
transform 1 0 -10898 0 1 5700
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_3
timestamp 1623563441
transform 1 0 6400 0 1 13720
box 0 2 400 98
use via_m1  via_m1_6
timestamp 1623561200
transform 1 0 -1698 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_2
timestamp 1623563441
transform 1 0 12000 0 1 13720
box 0 2 400 98
use via_m1  via_m1_7
timestamp 1623561200
transform 1 0 3902 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_1
timestamp 1623563441
transform 1 0 17600 0 1 13720
box 0 2 400 98
use via_m1  via_m1_10
timestamp 1623561200
transform 1 0 9502 0 1 6498
box 10898 6956 11298 7052
use via_m1  via_m1_11
timestamp 1623561200
transform 1 0 12302 0 1 5436
box 10898 6956 11298 7052
use power_ring  power_ring_0
timestamp 1623530672
transform 1 0 0 0 1 0
box 0 0 24400 21000
<< labels >>
flabel metal3 0 20600 5200 21000 1 FreeSans 16 0 0 0 vccd2
port 14 n power bidirectional
flabel metal3 18600 800 23600 1200 1 FreeSans 16 0 0 0 vssd2
port 15 s ground bidirectional
flabel metal2 13620 13898 13704 13982 1 FreeSans 16 0 0 0 p[8]
port 9 n signal output
flabel metal2 16748 13898 16832 13982 1 FreeSans 16 0 0 0 p[9]
port 10 nsew default output
flabel metal3 10308 13898 10392 13982 1 FreeSans 16 0 0 0 p[7]
port 8 n signal output
flabel metal2 5432 13898 5516 13982 1 FreeSans 16 0 0 0 p[6]
port 7 n signal output
flabel metal2 5062 7234 5146 7318 1 FreeSans 16 0 0 0 p[4]
port 5 s signal output
flabel metal2 8560 7234 8644 7318 1 FreeSans 16 0 0 0 p[3]
port 4 s signal output
flabel metal2 13160 7234 13244 7318 1 FreeSans 16 0 0 0 p[2]
port 3 s signal output
flabel metal2 15828 7234 15912 7318 1 FreeSans 16 0 0 0 p[1]
port 2 s signal output
flabel metal2 19232 7234 19316 7318 1 FreeSans 16 0 0 0 p[0]
port 1 s signal output
flabel metal2 1384 7234 1468 7318 1 FreeSans 16 0 0 0 p[5]
port 6 s signal output
flabel metal2 21164 13898 21248 13982 1 FreeSans 16 0 0 0 p[10]
port 11 n signal output
flabel metal2 24468 11442 24568 11542 1 FreeSans 16 0 0 0 input_analog
port 13 e signal input
flabel metal1 62 12378 142 12458 1 FreeSans 16 0 0 0 enb
port 12 w signal input
<< end >>
