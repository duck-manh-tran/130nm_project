magic
tech sky130A
timestamp 1623239895
<< pwell >>
rect -69 -105 536 605
<< nmos >>
rect 29 0 219 500
rect 248 0 438 500
<< ndiff >>
rect 0 483 29 500
rect 0 463 6 483
rect 23 463 29 483
rect 0 446 29 463
rect 0 426 6 446
rect 23 426 29 446
rect 0 409 29 426
rect 0 389 6 409
rect 23 389 29 409
rect 0 372 29 389
rect 0 352 6 372
rect 23 352 29 372
rect 0 335 29 352
rect 0 315 6 335
rect 23 315 29 335
rect 0 298 29 315
rect 0 278 6 298
rect 23 278 29 298
rect 0 261 29 278
rect 0 241 6 261
rect 23 241 29 261
rect 0 223 29 241
rect 0 203 6 223
rect 23 203 29 223
rect 0 186 29 203
rect 0 166 6 186
rect 23 166 29 186
rect 0 149 29 166
rect 0 129 6 149
rect 23 129 29 149
rect 0 112 29 129
rect 0 92 6 112
rect 23 92 29 112
rect 0 75 29 92
rect 0 55 6 75
rect 23 55 29 75
rect 0 38 29 55
rect 0 18 6 38
rect 23 18 29 38
rect 0 0 29 18
rect 219 483 248 500
rect 219 463 225 483
rect 242 463 248 483
rect 219 446 248 463
rect 219 426 225 446
rect 242 426 248 446
rect 219 409 248 426
rect 219 389 225 409
rect 242 389 248 409
rect 219 372 248 389
rect 219 352 225 372
rect 242 352 248 372
rect 219 335 248 352
rect 219 315 225 335
rect 242 315 248 335
rect 219 298 248 315
rect 219 278 225 298
rect 242 278 248 298
rect 219 261 248 278
rect 219 241 225 261
rect 242 241 248 261
rect 219 223 248 241
rect 219 203 225 223
rect 242 203 248 223
rect 219 186 248 203
rect 219 166 225 186
rect 242 166 248 186
rect 219 149 248 166
rect 219 129 225 149
rect 242 129 248 149
rect 219 112 248 129
rect 219 92 225 112
rect 242 92 248 112
rect 219 75 248 92
rect 219 55 225 75
rect 242 55 248 75
rect 219 38 248 55
rect 219 18 225 38
rect 242 18 248 38
rect 219 0 248 18
rect 438 483 467 500
rect 438 463 444 483
rect 461 463 467 483
rect 438 446 467 463
rect 438 426 444 446
rect 461 426 467 446
rect 438 409 467 426
rect 438 389 444 409
rect 461 389 467 409
rect 438 372 467 389
rect 438 352 444 372
rect 461 352 467 372
rect 438 335 467 352
rect 438 315 444 335
rect 461 315 467 335
rect 438 298 467 315
rect 438 278 444 298
rect 461 278 467 298
rect 438 261 467 278
rect 438 241 444 261
rect 461 241 467 261
rect 438 223 467 241
rect 438 203 444 223
rect 461 203 467 223
rect 438 186 467 203
rect 438 166 444 186
rect 461 166 467 186
rect 438 149 467 166
rect 438 129 444 149
rect 461 129 467 149
rect 438 112 467 129
rect 438 92 444 112
rect 461 92 467 112
rect 438 75 467 92
rect 438 55 444 75
rect 461 55 467 75
rect 438 38 467 55
rect 438 18 444 38
rect 461 18 467 38
rect 438 0 467 18
<< ndiffc >>
rect 6 463 23 483
rect 6 426 23 446
rect 6 389 23 409
rect 6 352 23 372
rect 6 315 23 335
rect 6 278 23 298
rect 6 241 23 261
rect 6 203 23 223
rect 6 166 23 186
rect 6 129 23 149
rect 6 92 23 112
rect 6 55 23 75
rect 6 18 23 38
rect 225 463 242 483
rect 225 426 242 446
rect 225 389 242 409
rect 225 352 242 372
rect 225 315 242 335
rect 225 278 242 298
rect 225 241 242 261
rect 225 203 242 223
rect 225 166 242 186
rect 225 129 242 149
rect 225 92 242 112
rect 225 55 242 75
rect 225 18 242 38
rect 444 463 461 483
rect 444 426 461 446
rect 444 389 461 409
rect 444 352 461 372
rect 444 315 461 335
rect 444 278 461 298
rect 444 241 461 261
rect 444 203 461 223
rect 444 166 461 186
rect 444 129 461 149
rect 444 92 461 112
rect 444 55 461 75
rect 444 18 461 38
<< poly >>
rect 29 500 219 544
rect 248 500 438 544
rect 29 -13 219 0
rect 248 -13 438 0
<< locali >>
rect 5 483 24 502
rect 5 463 6 483
rect 23 463 24 483
rect 5 446 24 463
rect 5 426 6 446
rect 23 426 24 446
rect 5 409 24 426
rect 5 389 6 409
rect 23 389 24 409
rect 5 372 24 389
rect 5 352 6 372
rect 23 352 24 372
rect 5 335 24 352
rect 5 315 6 335
rect 23 315 24 335
rect 5 298 24 315
rect 5 278 6 298
rect 23 278 24 298
rect 5 261 24 278
rect 5 241 6 261
rect 23 241 24 261
rect 5 223 24 241
rect 5 203 6 223
rect 23 203 24 223
rect 5 186 24 203
rect 5 166 6 186
rect 23 166 24 186
rect 5 149 24 166
rect 5 129 6 149
rect 23 129 24 149
rect 5 112 24 129
rect 5 92 6 112
rect 23 92 24 112
rect 5 75 24 92
rect 5 55 6 75
rect 23 55 24 75
rect 5 38 24 55
rect 5 18 6 38
rect 23 18 24 38
rect 5 -2 24 18
rect 224 483 243 502
rect 224 463 225 483
rect 242 463 243 483
rect 224 446 243 463
rect 224 426 225 446
rect 242 426 243 446
rect 224 409 243 426
rect 224 389 225 409
rect 242 389 243 409
rect 224 372 243 389
rect 224 352 225 372
rect 242 352 243 372
rect 224 335 243 352
rect 224 315 225 335
rect 242 315 243 335
rect 224 298 243 315
rect 224 278 225 298
rect 242 278 243 298
rect 224 261 243 278
rect 224 241 225 261
rect 242 241 243 261
rect 224 223 243 241
rect 224 203 225 223
rect 242 203 243 223
rect 224 186 243 203
rect 224 166 225 186
rect 242 166 243 186
rect 224 149 243 166
rect 224 129 225 149
rect 242 129 243 149
rect 224 112 243 129
rect 224 92 225 112
rect 242 92 243 112
rect 224 75 243 92
rect 224 55 225 75
rect 242 55 243 75
rect 224 38 243 55
rect 224 18 225 38
rect 242 18 243 38
rect 224 -2 243 18
rect 443 483 462 502
rect 443 463 444 483
rect 461 463 462 483
rect 443 446 462 463
rect 443 426 444 446
rect 461 426 462 446
rect 443 409 462 426
rect 443 389 444 409
rect 461 389 462 409
rect 443 372 462 389
rect 443 352 444 372
rect 461 352 462 372
rect 443 335 462 352
rect 443 315 444 335
rect 461 315 462 335
rect 443 298 462 315
rect 443 278 444 298
rect 461 278 462 298
rect 443 261 462 278
rect 443 241 444 261
rect 461 241 462 261
rect 443 223 462 241
rect 443 203 444 223
rect 461 203 462 223
rect 443 186 462 203
rect 443 166 444 186
rect 461 166 462 186
rect 443 149 462 166
rect 443 129 444 149
rect 461 129 462 149
rect 443 112 462 129
rect 443 92 444 112
rect 461 92 462 112
rect 443 75 462 92
rect 443 55 444 75
rect 461 55 462 75
rect 443 38 462 55
rect 443 18 444 38
rect 461 18 462 38
rect 443 -2 462 18
<< end >>
