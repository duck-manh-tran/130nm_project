magic
tech sky130A
magscale 1 2
timestamp 1623845735
<< ndiff >>
rect 1627 9858 1661 9892
<< pdiff >>
rect 1627 10182 1661 10216
<< locali >>
rect 1910 10148 1955 10192
rect 2308 10142 2353 10186
rect 1496 9984 1521 10018
<< metal1 >>
rect 0 10256 1994 10352
rect -90 9990 -10 10070
rect 21722 10004 23600 10076
rect 800 9712 1962 9808
<< metal2 >>
rect 5416 11416 5500 11500
rect 10290 11416 10374 11500
rect 13648 11416 13732 11500
rect 16708 11416 16792 11500
rect 21194 11416 21278 11500
rect 24520 9000 24620 9100
rect 1422 4856 1506 4940
rect 5050 4856 5134 4940
rect 8600 4856 8684 4940
rect 13198 4856 13282 4940
rect 15862 4856 15946 4940
rect 19222 4856 19306 4940
<< metal3 >>
rect 0 18200 5200 18600
rect 18600 -1600 23600 -1200
use via_m1  via_m1_4
timestamp 1623832439
transform 1 0 -7298 0 1 -1738
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_4
timestamp 1623832439
transform 1 0 6400 0 1 4960
box 0 2 400 98
use via_m1  via_m1_5
timestamp 1623832439
transform 1 0 -1698 0 1 -1738
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_5
timestamp 1623832439
transform 1 0 12000 0 1 4960
box 0 2 400 98
use via_m1  via_m1_8
timestamp 1623832439
transform 1 0 3902 0 1 -1738
box 10898 6956 11298 7052
use via_m1  via_m1_9
timestamp 1623832439
transform 1 0 9502 0 1 -1738
box 10898 6956 11298 7052
use via_m1  via_m1_3
timestamp 1623832439
transform 1 0 -7298 0 1 4098
box 10898 6956 11298 7052
use via_m1  via_m1_1
timestamp 1623832439
transform 1 0 -10898 0 1 3300
box 10898 6956 11298 7052
use via_m1  via_m1_2
timestamp 1623832439
transform 1 0 -10098 0 1 2756
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_3
timestamp 1623832439
transform 1 0 6400 0 1 11320
box 0 2 400 98
use via_m1  via_m1_6
timestamp 1623832439
transform 1 0 -1698 0 1 4098
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_2
timestamp 1623832439
transform 1 0 12000 0 1 11320
box 0 2 400 98
use via_m1  via_m1_7
timestamp 1623832439
transform 1 0 3902 0 1 4098
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_1
timestamp 1623832439
transform 1 0 17600 0 1 11320
box 0 2 400 98
use via_m1  via_m1_10
timestamp 1623832439
transform 1 0 9502 0 1 4098
box 10898 6956 11298 7052
use via_m1  via_m1_11
timestamp 1623832439
transform 1 0 12302 0 1 3036
box 10898 6956 11298 7052
use pwell_co_ring  pwell_co_ring_0
timestamp 1623832439
transform 1 0 3020 0 1 11340
box -1680 -6360 20145 60
use ring_osc  ring_osc_0
timestamp 1623845422
transform 1 0 1500 0 1 5200
box -1590 -344 23120 6300
use power_ring  power_ring_0
timestamp 1623832439
transform 1 0 0 0 1 -2400
box 0 0 24400 21000
<< labels >>
flabel metal1 -90 9990 -10 10070 1 FreeSans 16 0 0 0 enb
port 12 w signal input
flabel metal3 0 18200 5200 18600 1 FreeSans 16 0 0 0 vccd2
port 14 n power bidirectional
flabel metal3 18600 -1600 23600 -1200 1 FreeSans 16 0 0 0 vssd2
port 15 s ground bidirectional
flabel metal2 5416 11416 5500 11500 1 FreeSans 16 0 0 0 p[6]
port 7 n signal output
flabel metal2 10290 11416 10374 11500 1 FreeSans 16 0 0 0 p[7]
port 8 n signal output
flabel metal2 21194 11416 21278 11500 1 FreeSans 16 0 0 0 p[10]
port 11 n signal output
flabel metal2 19222 4856 19306 4940 1 FreeSans 16 0 0 0 p[0]
port 1 s signal output
flabel metal2 15862 4856 15946 4940 1 FreeSans 16 0 0 0 p[1]
port 2 s signal output
flabel metal2 13198 4856 13282 4940 1 FreeSans 16 0 0 0 p[2]
port 3 s signal output
flabel metal2 8600 4856 8684 4940 1 FreeSans 16 0 0 0 p[3]
port 4 s signal output
flabel metal2 5050 4856 5134 4940 1 FreeSans 16 0 0 0 p[4]
port 5 s signal output
flabel metal2 1422 4856 1506 4940 1 FreeSans 16 0 0 0 p[5]
port 6 s signal output
flabel metal2 16708 11416 16792 11500 1 FreeSans 16 0 0 0 p[9]
port 10 nsew default output
flabel metal2 24520 9000 24620 9100 1 FreeSans 16 0 0 0 input_analog
port 13 e signal input
flabel metal2 13648 11416 13732 11500 1 FreeSans 16 0 0 0 p[8]
port 9 n signal output
<< end >>
