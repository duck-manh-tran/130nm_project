VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO power_ring
  CLASS BLOCK ;
  FOREIGN power_ring ;
  ORIGIN 0.000 0.000 ;
  SIZE 122.000 BY 105.000 ;
  OBS
      LAYER met3 ;
        RECT 0.000 103.000 122.000 105.000 ;
        RECT 4.000 99.000 118.000 101.000 ;
        RECT 4.000 4.000 118.000 6.000 ;
        RECT 0.000 0.000 122.000 2.000 ;
      LAYER via3 ;
        RECT 0.200 104.400 0.600 104.800 ;
        RECT 0.800 104.400 1.200 104.800 ;
        RECT 1.400 104.400 1.800 104.800 ;
        RECT 18.200 104.400 18.600 104.800 ;
        RECT 18.800 104.400 19.200 104.800 ;
        RECT 19.400 104.400 19.800 104.800 ;
        RECT 46.200 104.400 46.600 104.800 ;
        RECT 46.800 104.400 47.200 104.800 ;
        RECT 47.400 104.400 47.800 104.800 ;
        RECT 74.200 104.400 74.600 104.800 ;
        RECT 74.800 104.400 75.200 104.800 ;
        RECT 75.400 104.400 75.800 104.800 ;
        RECT 102.200 104.400 102.600 104.800 ;
        RECT 102.800 104.400 103.200 104.800 ;
        RECT 103.400 104.400 103.800 104.800 ;
        RECT 120.200 104.400 120.600 104.800 ;
        RECT 120.800 104.400 121.200 104.800 ;
        RECT 121.400 104.400 121.800 104.800 ;
        RECT 0.200 103.800 0.600 104.200 ;
        RECT 0.800 103.800 1.200 104.200 ;
        RECT 1.400 103.800 1.800 104.200 ;
        RECT 18.200 103.800 18.600 104.200 ;
        RECT 18.800 103.800 19.200 104.200 ;
        RECT 19.400 103.800 19.800 104.200 ;
        RECT 46.200 103.800 46.600 104.200 ;
        RECT 46.800 103.800 47.200 104.200 ;
        RECT 47.400 103.800 47.800 104.200 ;
        RECT 74.200 103.800 74.600 104.200 ;
        RECT 74.800 103.800 75.200 104.200 ;
        RECT 75.400 103.800 75.800 104.200 ;
        RECT 102.200 103.800 102.600 104.200 ;
        RECT 102.800 103.800 103.200 104.200 ;
        RECT 103.400 103.800 103.800 104.200 ;
        RECT 120.200 103.800 120.600 104.200 ;
        RECT 120.800 103.800 121.200 104.200 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 0.200 103.200 0.600 103.600 ;
        RECT 0.800 103.200 1.200 103.600 ;
        RECT 1.400 103.200 1.800 103.600 ;
        RECT 18.200 103.200 18.600 103.600 ;
        RECT 18.800 103.200 19.200 103.600 ;
        RECT 19.400 103.200 19.800 103.600 ;
        RECT 46.200 103.200 46.600 103.600 ;
        RECT 46.800 103.200 47.200 103.600 ;
        RECT 47.400 103.200 47.800 103.600 ;
        RECT 74.200 103.200 74.600 103.600 ;
        RECT 74.800 103.200 75.200 103.600 ;
        RECT 75.400 103.200 75.800 103.600 ;
        RECT 102.200 103.200 102.600 103.600 ;
        RECT 102.800 103.200 103.200 103.600 ;
        RECT 103.400 103.200 103.800 103.600 ;
        RECT 120.200 103.200 120.600 103.600 ;
        RECT 120.800 103.200 121.200 103.600 ;
        RECT 121.400 103.200 121.800 103.600 ;
        RECT 4.200 100.400 4.600 100.800 ;
        RECT 4.800 100.400 5.200 100.800 ;
        RECT 5.400 100.400 5.800 100.800 ;
        RECT 32.200 100.400 32.600 100.800 ;
        RECT 32.800 100.400 33.200 100.800 ;
        RECT 33.400 100.400 33.800 100.800 ;
        RECT 60.200 100.400 60.600 100.800 ;
        RECT 60.800 100.400 61.200 100.800 ;
        RECT 61.400 100.400 61.800 100.800 ;
        RECT 88.200 100.400 88.600 100.800 ;
        RECT 88.800 100.400 89.200 100.800 ;
        RECT 89.400 100.400 89.800 100.800 ;
        RECT 116.200 100.400 116.600 100.800 ;
        RECT 116.800 100.400 117.200 100.800 ;
        RECT 117.400 100.400 117.800 100.800 ;
        RECT 4.200 99.800 4.600 100.200 ;
        RECT 4.800 99.800 5.200 100.200 ;
        RECT 5.400 99.800 5.800 100.200 ;
        RECT 32.200 99.800 32.600 100.200 ;
        RECT 32.800 99.800 33.200 100.200 ;
        RECT 33.400 99.800 33.800 100.200 ;
        RECT 60.200 99.800 60.600 100.200 ;
        RECT 60.800 99.800 61.200 100.200 ;
        RECT 61.400 99.800 61.800 100.200 ;
        RECT 88.200 99.800 88.600 100.200 ;
        RECT 88.800 99.800 89.200 100.200 ;
        RECT 89.400 99.800 89.800 100.200 ;
        RECT 116.200 99.800 116.600 100.200 ;
        RECT 116.800 99.800 117.200 100.200 ;
        RECT 117.400 99.800 117.800 100.200 ;
        RECT 4.200 99.200 4.600 99.600 ;
        RECT 4.800 99.200 5.200 99.600 ;
        RECT 5.400 99.200 5.800 99.600 ;
        RECT 32.200 99.200 32.600 99.600 ;
        RECT 32.800 99.200 33.200 99.600 ;
        RECT 33.400 99.200 33.800 99.600 ;
        RECT 60.200 99.200 60.600 99.600 ;
        RECT 60.800 99.200 61.200 99.600 ;
        RECT 61.400 99.200 61.800 99.600 ;
        RECT 88.200 99.200 88.600 99.600 ;
        RECT 88.800 99.200 89.200 99.600 ;
        RECT 89.400 99.200 89.800 99.600 ;
        RECT 116.200 99.200 116.600 99.600 ;
        RECT 116.800 99.200 117.200 99.600 ;
        RECT 117.400 99.200 117.800 99.600 ;
        RECT 4.200 5.400 4.600 5.800 ;
        RECT 4.800 5.400 5.200 5.800 ;
        RECT 5.400 5.400 5.800 5.800 ;
        RECT 32.200 5.400 32.600 5.800 ;
        RECT 32.800 5.400 33.200 5.800 ;
        RECT 33.400 5.400 33.800 5.800 ;
        RECT 60.200 5.400 60.600 5.800 ;
        RECT 60.800 5.400 61.200 5.800 ;
        RECT 61.400 5.400 61.800 5.800 ;
        RECT 88.200 5.400 88.600 5.800 ;
        RECT 88.800 5.400 89.200 5.800 ;
        RECT 89.400 5.400 89.800 5.800 ;
        RECT 116.200 5.400 116.600 5.800 ;
        RECT 116.800 5.400 117.200 5.800 ;
        RECT 117.400 5.400 117.800 5.800 ;
        RECT 4.200 4.800 4.600 5.200 ;
        RECT 4.800 4.800 5.200 5.200 ;
        RECT 5.400 4.800 5.800 5.200 ;
        RECT 32.200 4.800 32.600 5.200 ;
        RECT 32.800 4.800 33.200 5.200 ;
        RECT 33.400 4.800 33.800 5.200 ;
        RECT 60.200 4.800 60.600 5.200 ;
        RECT 60.800 4.800 61.200 5.200 ;
        RECT 61.400 4.800 61.800 5.200 ;
        RECT 88.200 4.800 88.600 5.200 ;
        RECT 88.800 4.800 89.200 5.200 ;
        RECT 89.400 4.800 89.800 5.200 ;
        RECT 116.200 4.800 116.600 5.200 ;
        RECT 116.800 4.800 117.200 5.200 ;
        RECT 117.400 4.800 117.800 5.200 ;
        RECT 4.200 4.200 4.600 4.600 ;
        RECT 4.800 4.200 5.200 4.600 ;
        RECT 5.400 4.200 5.800 4.600 ;
        RECT 32.200 4.200 32.600 4.600 ;
        RECT 32.800 4.200 33.200 4.600 ;
        RECT 33.400 4.200 33.800 4.600 ;
        RECT 60.200 4.200 60.600 4.600 ;
        RECT 60.800 4.200 61.200 4.600 ;
        RECT 61.400 4.200 61.800 4.600 ;
        RECT 88.200 4.200 88.600 4.600 ;
        RECT 88.800 4.200 89.200 4.600 ;
        RECT 89.400 4.200 89.800 4.600 ;
        RECT 116.200 4.200 116.600 4.600 ;
        RECT 116.800 4.200 117.200 4.600 ;
        RECT 117.400 4.200 117.800 4.600 ;
        RECT 0.200 1.400 0.600 1.800 ;
        RECT 0.800 1.400 1.200 1.800 ;
        RECT 1.400 1.400 1.800 1.800 ;
        RECT 18.200 1.400 18.600 1.800 ;
        RECT 18.800 1.400 19.200 1.800 ;
        RECT 19.400 1.400 19.800 1.800 ;
        RECT 46.200 1.400 46.600 1.800 ;
        RECT 46.800 1.400 47.200 1.800 ;
        RECT 47.400 1.400 47.800 1.800 ;
        RECT 74.200 1.400 74.600 1.800 ;
        RECT 74.800 1.400 75.200 1.800 ;
        RECT 75.400 1.400 75.800 1.800 ;
        RECT 102.200 1.400 102.600 1.800 ;
        RECT 102.800 1.400 103.200 1.800 ;
        RECT 103.400 1.400 103.800 1.800 ;
        RECT 120.200 1.400 120.600 1.800 ;
        RECT 120.800 1.400 121.200 1.800 ;
        RECT 121.400 1.400 121.800 1.800 ;
        RECT 0.200 0.800 0.600 1.200 ;
        RECT 0.800 0.800 1.200 1.200 ;
        RECT 1.400 0.800 1.800 1.200 ;
        RECT 18.200 0.800 18.600 1.200 ;
        RECT 18.800 0.800 19.200 1.200 ;
        RECT 19.400 0.800 19.800 1.200 ;
        RECT 46.200 0.800 46.600 1.200 ;
        RECT 46.800 0.800 47.200 1.200 ;
        RECT 47.400 0.800 47.800 1.200 ;
        RECT 74.200 0.800 74.600 1.200 ;
        RECT 74.800 0.800 75.200 1.200 ;
        RECT 75.400 0.800 75.800 1.200 ;
        RECT 102.200 0.800 102.600 1.200 ;
        RECT 102.800 0.800 103.200 1.200 ;
        RECT 103.400 0.800 103.800 1.200 ;
        RECT 120.200 0.800 120.600 1.200 ;
        RECT 120.800 0.800 121.200 1.200 ;
        RECT 121.400 0.800 121.800 1.200 ;
        RECT 0.200 0.200 0.600 0.600 ;
        RECT 0.800 0.200 1.200 0.600 ;
        RECT 1.400 0.200 1.800 0.600 ;
        RECT 18.200 0.200 18.600 0.600 ;
        RECT 18.800 0.200 19.200 0.600 ;
        RECT 19.400 0.200 19.800 0.600 ;
        RECT 46.200 0.200 46.600 0.600 ;
        RECT 46.800 0.200 47.200 0.600 ;
        RECT 47.400 0.200 47.800 0.600 ;
        RECT 74.200 0.200 74.600 0.600 ;
        RECT 74.800 0.200 75.200 0.600 ;
        RECT 75.400 0.200 75.800 0.600 ;
        RECT 102.200 0.200 102.600 0.600 ;
        RECT 102.800 0.200 103.200 0.600 ;
        RECT 103.400 0.200 103.800 0.600 ;
        RECT 120.200 0.200 120.600 0.600 ;
        RECT 120.800 0.200 121.200 0.600 ;
        RECT 121.400 0.200 121.800 0.600 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 105.000 ;
        RECT 4.000 4.000 6.000 101.000 ;
        RECT 18.000 0.000 20.000 105.000 ;
        RECT 32.000 4.000 34.000 101.000 ;
        RECT 46.000 0.000 48.000 105.000 ;
        RECT 60.000 4.000 62.000 101.000 ;
        RECT 74.000 0.000 76.000 105.000 ;
        RECT 88.000 4.000 90.000 101.000 ;
        RECT 102.000 0.000 104.000 105.000 ;
        RECT 116.000 4.000 118.000 101.000 ;
        RECT 120.000 0.000 122.000 105.000 ;
  END
END power_ring
MACRO pwell_co_ring
  CLASS BLOCK ;
  FOREIGN pwell_co_ring ;
  ORIGIN 8.400 31.800 ;
  SIZE 109.125 BY 32.100 ;
  OBS
      LAYER li1 ;
        RECT -0.100 0.000 90.900 0.300 ;
        RECT -0.100 -15.630 0.200 0.000 ;
        RECT 90.600 -15.630 90.900 0.000 ;
        RECT -8.400 -15.930 100.725 -15.630 ;
        RECT -8.400 -31.500 -8.100 -15.930 ;
        RECT 100.400 -16.000 100.725 -15.930 ;
        RECT 100.400 -31.500 100.700 -16.000 ;
        RECT -8.400 -31.800 100.700 -31.500 ;
  END
END pwell_co_ring
MACRO via_m4_li
  CLASS BLOCK ;
  FOREIGN via_m4_li ;
  ORIGIN 0.000 -0.010 ;
  SIZE 2.000 BY 0.480 ;
  OBS
      LAYER li1 ;
        RECT 0.000 0.100 2.000 0.400 ;
      LAYER mcon ;
        RECT 0.110 0.100 0.410 0.400 ;
        RECT 0.600 0.100 0.900 0.400 ;
        RECT 1.100 0.100 1.400 0.400 ;
        RECT 1.590 0.100 1.890 0.400 ;
      LAYER met1 ;
        RECT 0.080 0.010 1.920 0.490 ;
      LAYER via ;
        RECT 0.130 0.100 0.430 0.400 ;
        RECT 0.490 0.100 0.790 0.400 ;
        RECT 0.850 0.100 1.150 0.400 ;
        RECT 1.210 0.100 1.510 0.400 ;
        RECT 1.570 0.100 1.870 0.400 ;
      LAYER met2 ;
        RECT 0.000 0.010 2.000 0.490 ;
      LAYER via2 ;
        RECT 0.180 0.090 0.500 0.410 ;
        RECT 0.620 0.090 0.940 0.410 ;
        RECT 1.060 0.090 1.380 0.410 ;
        RECT 1.500 0.090 1.820 0.410 ;
      LAYER met3 ;
        RECT 0.000 0.010 2.000 0.490 ;
      LAYER via3 ;
        RECT 0.160 0.070 0.520 0.435 ;
        RECT 0.600 0.070 0.960 0.435 ;
        RECT 1.040 0.070 1.400 0.435 ;
        RECT 1.480 0.070 1.840 0.435 ;
      LAYER met4 ;
        RECT 0.000 0.010 2.000 0.490 ;
  END
END via_m4_li
MACRO via_m1
  CLASS BLOCK ;
  FOREIGN via_m1 ;
  ORIGIN -54.490 -34.780 ;
  SIZE 2.000 BY 0.480 ;
  OBS
      LAYER met1 ;
        RECT 54.620 34.780 56.360 35.260 ;
      LAYER via ;
        RECT 54.620 34.870 54.920 35.170 ;
        RECT 54.980 34.870 55.280 35.170 ;
        RECT 55.340 34.870 55.640 35.170 ;
        RECT 55.700 34.870 56.000 35.170 ;
        RECT 56.060 34.870 56.360 35.170 ;
      LAYER met2 ;
        RECT 54.490 34.780 56.490 35.260 ;
      LAYER via2 ;
        RECT 54.670 34.860 54.990 35.180 ;
        RECT 55.110 34.860 55.430 35.180 ;
        RECT 55.550 34.860 55.870 35.180 ;
        RECT 55.990 34.860 56.310 35.180 ;
      LAYER met3 ;
        RECT 54.490 34.780 56.490 35.260 ;
      LAYER via3 ;
        RECT 54.650 34.840 55.010 35.205 ;
        RECT 55.090 34.840 55.450 35.205 ;
        RECT 55.530 34.840 55.890 35.205 ;
        RECT 55.970 34.840 56.330 35.205 ;
      LAYER met4 ;
        RECT 54.490 34.780 56.490 35.260 ;
  END
END via_m1
MACRO ring_osc
  CLASS BLOCK ;
  FOREIGN ring_osc ;
  ORIGIN 2.510 0.000 ;
  SIZE 111.870 BY 29.840 ;
  OBS
      LAYER nwell ;
        RECT -1.000 24.105 1.680 25.950 ;
        RECT 2.995 24.105 4.755 25.710 ;
      LAYER pwell ;
        RECT -0.320 23.585 1.485 23.815 ;
        RECT -0.805 22.905 1.485 23.585 ;
      LAYER nwell ;
        RECT 8.480 22.965 97.550 29.840 ;
        RECT 19.520 22.960 26.710 22.965 ;
        RECT 37.230 22.960 44.420 22.965 ;
        RECT 54.940 22.960 62.130 22.965 ;
        RECT 72.650 22.960 79.840 22.965 ;
        RECT 90.360 22.960 97.550 22.965 ;
      LAYER pwell ;
        RECT -0.660 22.715 -0.490 22.905 ;
        RECT 3.330 22.715 3.500 22.885 ;
        RECT 8.480 15.470 97.550 22.570 ;
        RECT 100.500 20.000 103.500 25.000 ;
        RECT 100.500 19.000 108.500 20.000 ;
        RECT 102.500 17.000 108.500 19.000 ;
        RECT 0.000 7.270 106.780 14.370 ;
      LAYER nwell ;
        RECT 0.000 6.875 7.190 6.880 ;
        RECT 17.710 6.875 24.900 6.880 ;
        RECT 35.420 6.875 42.610 6.880 ;
        RECT 53.130 6.875 60.320 6.880 ;
        RECT 70.840 6.875 78.030 6.880 ;
        RECT 88.550 6.875 95.740 6.880 ;
        RECT 0.000 0.000 106.780 6.875 ;
      LAYER li1 ;
        RECT 8.660 29.660 10.550 29.690 ;
        RECT 12.340 29.660 16.190 29.690 ;
        RECT 17.850 29.660 21.700 29.690 ;
        RECT 23.540 29.660 24.940 29.690 ;
        RECT 26.370 29.660 28.260 29.690 ;
        RECT 30.050 29.660 33.900 29.690 ;
        RECT 35.560 29.660 39.410 29.690 ;
        RECT 41.250 29.660 42.650 29.690 ;
        RECT 44.080 29.660 45.970 29.690 ;
        RECT 47.760 29.660 51.610 29.690 ;
        RECT 53.270 29.660 57.120 29.690 ;
        RECT 58.960 29.660 60.360 29.690 ;
        RECT 61.790 29.660 63.680 29.690 ;
        RECT 65.470 29.660 69.320 29.690 ;
        RECT 70.980 29.660 74.830 29.690 ;
        RECT 76.670 29.660 78.070 29.690 ;
        RECT 79.500 29.660 81.390 29.690 ;
        RECT 83.180 29.660 87.030 29.690 ;
        RECT 88.690 29.660 92.540 29.690 ;
        RECT 94.380 29.660 95.780 29.690 ;
        RECT 8.660 29.490 97.370 29.660 ;
        RECT 8.660 29.330 10.550 29.490 ;
        RECT 12.340 29.330 16.190 29.490 ;
        RECT 17.850 29.330 21.700 29.490 ;
        RECT 23.540 29.330 24.940 29.490 ;
        RECT 26.370 29.330 28.260 29.490 ;
        RECT 30.050 29.330 33.900 29.490 ;
        RECT 35.560 29.330 39.410 29.490 ;
        RECT 41.250 29.330 42.650 29.490 ;
        RECT 44.080 29.330 45.970 29.490 ;
        RECT 47.760 29.330 51.610 29.490 ;
        RECT 53.270 29.330 57.120 29.490 ;
        RECT 58.960 29.330 60.360 29.490 ;
        RECT 61.790 29.330 63.680 29.490 ;
        RECT 65.470 29.330 69.320 29.490 ;
        RECT 70.980 29.330 74.830 29.490 ;
        RECT 76.670 29.330 78.070 29.490 ;
        RECT 79.500 29.330 81.390 29.490 ;
        RECT 83.180 29.330 87.030 29.490 ;
        RECT 88.690 29.330 92.540 29.490 ;
        RECT 94.380 29.330 95.780 29.490 ;
        RECT -0.810 25.605 0.190 25.770 ;
        RECT -0.810 25.435 1.490 25.605 ;
        RECT 3.185 25.435 4.565 25.605 ;
        RECT -0.725 24.865 -0.465 25.265 ;
        RECT -0.295 25.035 0.640 25.435 ;
        RECT 0.810 24.925 1.405 25.265 ;
        RECT -0.725 24.695 0.640 24.865 ;
        RECT -0.725 23.795 -0.265 24.525 ;
        RECT -0.095 23.625 0.640 24.695 ;
        RECT -0.725 23.455 0.640 23.625 ;
        RECT 0.810 23.605 0.985 24.925 ;
        RECT 1.165 24.750 1.405 24.755 ;
        RECT 1.680 24.750 3.005 24.960 ;
        RECT 1.165 24.740 3.005 24.750 ;
        RECT 1.165 24.530 1.900 24.740 ;
        RECT 2.785 24.535 3.005 24.740 ;
        RECT 3.460 24.710 3.790 25.435 ;
        RECT 3.270 24.535 3.790 24.540 ;
        RECT 1.165 23.775 1.405 24.530 ;
        RECT 2.785 24.315 3.790 24.535 ;
        RECT 0.810 23.480 1.405 23.605 ;
        RECT 2.210 23.480 2.510 24.310 ;
        RECT -0.725 23.055 -0.465 23.455 ;
        RECT -0.295 22.885 0.640 23.285 ;
        RECT 0.810 23.180 2.510 23.480 ;
        RECT 0.810 23.055 1.405 23.180 ;
        RECT 3.270 23.055 3.790 24.315 ;
        RECT 3.960 23.715 4.480 25.265 ;
        RECT 8.660 24.460 8.830 29.330 ;
        RECT 9.170 24.040 9.460 29.330 ;
        RECT 3.960 22.885 4.300 23.545 ;
        RECT 10.380 22.950 10.760 23.000 ;
        RECT -0.810 22.715 1.490 22.885 ;
        RECT 3.185 22.715 4.565 22.885 ;
        RECT 9.430 22.590 10.760 22.950 ;
        RECT 10.380 22.540 10.760 22.590 ;
        RECT 9.170 16.090 9.460 21.540 ;
        RECT 11.355 16.500 11.655 29.090 ;
        RECT 13.550 24.040 13.840 29.330 ;
        RECT 14.180 24.460 14.350 29.330 ;
        RECT 14.690 24.040 14.980 29.330 ;
        RECT 12.250 22.950 12.630 23.000 ;
        RECT 15.900 22.950 16.280 23.000 ;
        RECT 12.250 22.590 13.580 22.950 ;
        RECT 14.950 22.590 16.280 22.950 ;
        RECT 12.250 22.540 12.630 22.590 ;
        RECT 15.900 22.540 16.280 22.590 ;
        RECT 13.550 16.090 13.840 21.540 ;
        RECT 14.690 16.090 14.980 21.540 ;
        RECT 16.875 16.500 17.175 29.090 ;
        RECT 19.070 24.040 19.360 29.330 ;
        RECT 19.700 24.460 19.870 29.330 ;
        RECT 20.210 24.030 20.500 29.330 ;
        RECT 17.770 22.950 18.150 23.000 ;
        RECT 21.420 22.950 21.800 23.000 ;
        RECT 17.770 22.590 19.100 22.950 ;
        RECT 20.470 22.590 21.800 22.950 ;
        RECT 17.770 22.540 18.150 22.590 ;
        RECT 21.420 22.540 21.800 22.590 ;
        RECT 19.070 16.090 19.360 21.540 ;
        RECT 20.210 16.090 20.500 21.540 ;
        RECT 22.400 16.500 22.700 29.090 ;
        RECT 23.540 24.030 23.830 29.330 ;
        RECT 24.750 22.950 25.130 23.000 ;
        RECT 23.800 22.590 25.130 22.950 ;
        RECT 24.750 22.540 25.130 22.590 ;
        RECT 23.540 16.090 23.830 21.540 ;
        RECT 25.730 16.500 26.030 29.090 ;
        RECT 26.370 24.460 26.540 29.330 ;
        RECT 26.880 24.040 27.170 29.330 ;
        RECT 28.090 22.950 28.470 23.000 ;
        RECT 27.140 22.590 28.470 22.950 ;
        RECT 28.090 22.540 28.470 22.590 ;
        RECT 26.880 16.090 27.170 21.540 ;
        RECT 29.065 16.500 29.365 29.090 ;
        RECT 31.260 24.040 31.550 29.330 ;
        RECT 31.890 24.460 32.060 29.330 ;
        RECT 32.400 24.040 32.690 29.330 ;
        RECT 29.960 22.950 30.340 23.000 ;
        RECT 33.610 22.950 33.990 23.000 ;
        RECT 29.960 22.590 31.290 22.950 ;
        RECT 32.660 22.590 33.990 22.950 ;
        RECT 29.960 22.540 30.340 22.590 ;
        RECT 33.610 22.540 33.990 22.590 ;
        RECT 31.260 16.090 31.550 21.540 ;
        RECT 32.400 16.090 32.690 21.540 ;
        RECT 34.585 16.500 34.885 29.090 ;
        RECT 36.780 24.040 37.070 29.330 ;
        RECT 37.410 24.460 37.580 29.330 ;
        RECT 37.920 24.030 38.210 29.330 ;
        RECT 35.480 22.950 35.860 23.000 ;
        RECT 39.130 22.950 39.510 23.000 ;
        RECT 35.480 22.590 36.810 22.950 ;
        RECT 38.180 22.590 39.510 22.950 ;
        RECT 35.480 22.540 35.860 22.590 ;
        RECT 39.130 22.540 39.510 22.590 ;
        RECT 36.780 16.090 37.070 21.540 ;
        RECT 37.920 16.090 38.210 21.540 ;
        RECT 40.110 16.500 40.410 29.090 ;
        RECT 41.250 24.030 41.540 29.330 ;
        RECT 42.460 22.950 42.840 23.000 ;
        RECT 41.510 22.590 42.840 22.950 ;
        RECT 42.460 22.540 42.840 22.590 ;
        RECT 41.250 16.090 41.540 21.540 ;
        RECT 43.440 16.500 43.740 29.090 ;
        RECT 44.080 24.460 44.250 29.330 ;
        RECT 44.590 24.040 44.880 29.330 ;
        RECT 45.800 22.950 46.180 23.000 ;
        RECT 44.850 22.590 46.180 22.950 ;
        RECT 45.800 22.540 46.180 22.590 ;
        RECT 44.590 16.090 44.880 21.540 ;
        RECT 46.775 16.500 47.075 29.090 ;
        RECT 48.970 24.040 49.260 29.330 ;
        RECT 49.600 24.460 49.770 29.330 ;
        RECT 50.110 24.040 50.400 29.330 ;
        RECT 47.670 22.950 48.050 23.000 ;
        RECT 51.320 22.950 51.700 23.000 ;
        RECT 47.670 22.590 49.000 22.950 ;
        RECT 50.370 22.590 51.700 22.950 ;
        RECT 47.670 22.540 48.050 22.590 ;
        RECT 51.320 22.540 51.700 22.590 ;
        RECT 48.970 16.090 49.260 21.540 ;
        RECT 50.110 16.090 50.400 21.540 ;
        RECT 52.295 16.500 52.595 29.090 ;
        RECT 54.490 24.040 54.780 29.330 ;
        RECT 55.120 24.460 55.290 29.330 ;
        RECT 55.630 24.030 55.920 29.330 ;
        RECT 53.190 22.950 53.570 23.000 ;
        RECT 56.840 22.950 57.220 23.000 ;
        RECT 53.190 22.590 54.520 22.950 ;
        RECT 55.890 22.590 57.220 22.950 ;
        RECT 53.190 22.540 53.570 22.590 ;
        RECT 56.840 22.540 57.220 22.590 ;
        RECT 54.490 16.090 54.780 21.540 ;
        RECT 55.630 16.090 55.920 21.540 ;
        RECT 57.820 16.500 58.120 29.090 ;
        RECT 58.960 24.030 59.250 29.330 ;
        RECT 60.170 22.950 60.550 23.000 ;
        RECT 59.220 22.590 60.550 22.950 ;
        RECT 60.170 22.540 60.550 22.590 ;
        RECT 58.960 16.090 59.250 21.540 ;
        RECT 61.150 16.500 61.450 29.090 ;
        RECT 61.790 24.460 61.960 29.330 ;
        RECT 62.300 24.040 62.590 29.330 ;
        RECT 63.510 22.950 63.890 23.000 ;
        RECT 62.560 22.590 63.890 22.950 ;
        RECT 63.510 22.540 63.890 22.590 ;
        RECT 62.300 16.090 62.590 21.540 ;
        RECT 64.485 16.500 64.785 29.090 ;
        RECT 66.680 24.040 66.970 29.330 ;
        RECT 67.310 24.460 67.480 29.330 ;
        RECT 67.820 24.040 68.110 29.330 ;
        RECT 65.380 22.950 65.760 23.000 ;
        RECT 69.030 22.950 69.410 23.000 ;
        RECT 65.380 22.590 66.710 22.950 ;
        RECT 68.080 22.590 69.410 22.950 ;
        RECT 65.380 22.540 65.760 22.590 ;
        RECT 69.030 22.540 69.410 22.590 ;
        RECT 66.680 16.090 66.970 21.540 ;
        RECT 67.820 16.090 68.110 21.540 ;
        RECT 70.005 16.500 70.305 29.090 ;
        RECT 72.200 24.040 72.490 29.330 ;
        RECT 72.830 24.460 73.000 29.330 ;
        RECT 73.340 24.030 73.630 29.330 ;
        RECT 70.900 22.950 71.280 23.000 ;
        RECT 74.550 22.950 74.930 23.000 ;
        RECT 70.900 22.590 72.230 22.950 ;
        RECT 73.600 22.590 74.930 22.950 ;
        RECT 70.900 22.540 71.280 22.590 ;
        RECT 74.550 22.540 74.930 22.590 ;
        RECT 72.200 16.090 72.490 21.540 ;
        RECT 73.340 16.090 73.630 21.540 ;
        RECT 75.530 16.500 75.830 29.090 ;
        RECT 76.670 24.030 76.960 29.330 ;
        RECT 77.880 22.950 78.260 23.000 ;
        RECT 76.930 22.590 78.260 22.950 ;
        RECT 77.880 22.540 78.260 22.590 ;
        RECT 76.670 16.090 76.960 21.540 ;
        RECT 78.860 16.500 79.160 29.090 ;
        RECT 79.500 24.460 79.670 29.330 ;
        RECT 80.010 24.040 80.300 29.330 ;
        RECT 81.220 22.950 81.600 23.000 ;
        RECT 80.270 22.590 81.600 22.950 ;
        RECT 81.220 22.540 81.600 22.590 ;
        RECT 80.010 16.090 80.300 21.540 ;
        RECT 82.195 16.500 82.495 29.090 ;
        RECT 84.390 24.040 84.680 29.330 ;
        RECT 85.020 24.460 85.190 29.330 ;
        RECT 85.530 24.040 85.820 29.330 ;
        RECT 83.090 22.950 83.470 23.000 ;
        RECT 86.740 22.950 87.120 23.000 ;
        RECT 83.090 22.590 84.420 22.950 ;
        RECT 85.790 22.590 87.120 22.950 ;
        RECT 83.090 22.540 83.470 22.590 ;
        RECT 86.740 22.540 87.120 22.590 ;
        RECT 84.390 16.090 84.680 21.540 ;
        RECT 85.530 16.090 85.820 21.540 ;
        RECT 87.715 16.500 88.015 29.090 ;
        RECT 89.910 24.040 90.200 29.330 ;
        RECT 90.540 24.460 90.710 29.330 ;
        RECT 91.050 24.030 91.340 29.330 ;
        RECT 88.610 22.950 88.990 23.000 ;
        RECT 92.260 22.950 92.640 23.000 ;
        RECT 88.610 22.590 89.940 22.950 ;
        RECT 91.310 22.590 92.640 22.950 ;
        RECT 88.610 22.540 88.990 22.590 ;
        RECT 92.260 22.540 92.640 22.590 ;
        RECT 89.910 16.090 90.200 21.540 ;
        RECT 91.050 16.090 91.340 21.540 ;
        RECT 93.240 16.500 93.540 29.090 ;
        RECT 94.380 24.030 94.670 29.330 ;
        RECT 95.590 22.950 95.970 23.000 ;
        RECT 94.640 22.590 95.970 22.950 ;
        RECT 95.590 22.540 95.970 22.590 ;
        RECT 94.380 16.090 94.670 21.540 ;
        RECT 96.570 16.500 96.870 29.090 ;
        RECT 101.000 24.015 103.000 24.380 ;
        RECT 101.000 19.500 103.000 19.865 ;
        RECT 102.000 18.500 103.365 19.500 ;
        RECT 103.000 17.500 103.365 18.500 ;
        RECT 107.515 18.500 108.500 19.500 ;
        RECT 107.515 17.500 107.880 18.500 ;
        RECT 8.660 15.730 10.550 16.090 ;
        RECT 12.340 15.730 16.190 16.090 ;
        RECT 17.850 15.730 21.700 16.090 ;
        RECT 23.540 15.730 24.940 16.090 ;
        RECT 26.370 15.730 28.260 16.090 ;
        RECT 30.050 15.730 33.900 16.090 ;
        RECT 35.560 15.730 39.410 16.090 ;
        RECT 41.250 15.730 42.650 16.090 ;
        RECT 44.080 15.730 45.970 16.090 ;
        RECT 47.760 15.730 51.610 16.090 ;
        RECT 53.270 15.730 57.120 16.090 ;
        RECT 58.960 15.730 60.360 16.090 ;
        RECT 61.790 15.730 63.680 16.090 ;
        RECT 65.470 15.730 69.320 16.090 ;
        RECT 70.980 15.730 74.830 16.090 ;
        RECT 76.670 15.730 78.070 16.090 ;
        RECT 79.500 15.730 81.390 16.090 ;
        RECT 83.180 15.730 87.030 16.090 ;
        RECT 88.690 15.730 92.540 16.090 ;
        RECT 94.380 15.730 95.780 16.090 ;
        RECT 1.770 13.750 3.170 14.110 ;
        RECT 5.010 13.750 8.860 14.110 ;
        RECT 10.520 13.750 14.370 14.110 ;
        RECT 16.160 13.750 18.050 14.110 ;
        RECT 19.480 13.750 20.880 14.110 ;
        RECT 22.720 13.750 26.570 14.110 ;
        RECT 28.230 13.750 32.080 14.110 ;
        RECT 33.870 13.750 35.760 14.110 ;
        RECT 37.190 13.750 38.590 14.110 ;
        RECT 40.430 13.750 44.280 14.110 ;
        RECT 45.940 13.750 49.790 14.110 ;
        RECT 51.580 13.750 53.470 14.110 ;
        RECT 54.900 13.750 56.300 14.110 ;
        RECT 58.140 13.750 61.990 14.110 ;
        RECT 63.650 13.750 67.500 14.110 ;
        RECT 69.290 13.750 71.180 14.110 ;
        RECT 72.610 13.750 74.010 14.110 ;
        RECT 75.850 13.750 79.700 14.110 ;
        RECT 81.360 13.750 85.210 14.110 ;
        RECT 87.000 13.750 88.890 14.110 ;
        RECT 90.320 13.750 91.720 14.110 ;
        RECT 93.560 13.750 97.410 14.110 ;
        RECT 99.070 13.750 102.920 14.110 ;
        RECT 104.710 13.750 106.600 14.110 ;
        RECT 0.680 0.750 0.980 13.340 ;
        RECT 2.880 8.300 3.170 13.750 ;
        RECT 1.580 7.250 1.960 7.300 ;
        RECT 1.580 6.890 2.910 7.250 ;
        RECT 1.580 6.840 1.960 6.890 ;
        RECT 2.880 0.510 3.170 5.810 ;
        RECT 4.010 0.750 4.310 13.340 ;
        RECT 6.210 8.300 6.500 13.750 ;
        RECT 7.350 8.300 7.640 13.750 ;
        RECT 4.910 7.250 5.290 7.300 ;
        RECT 8.560 7.250 8.940 7.300 ;
        RECT 4.910 6.890 6.240 7.250 ;
        RECT 7.610 6.890 8.940 7.250 ;
        RECT 4.910 6.840 5.290 6.890 ;
        RECT 8.560 6.840 8.940 6.890 ;
        RECT 6.210 0.510 6.500 5.810 ;
        RECT 6.840 0.510 7.010 5.380 ;
        RECT 7.350 0.510 7.640 5.800 ;
        RECT 9.535 0.750 9.835 13.340 ;
        RECT 11.730 8.300 12.020 13.750 ;
        RECT 12.870 8.300 13.160 13.750 ;
        RECT 10.430 7.250 10.810 7.300 ;
        RECT 14.080 7.250 14.460 7.300 ;
        RECT 10.430 6.890 11.760 7.250 ;
        RECT 13.130 6.890 14.460 7.250 ;
        RECT 10.430 6.840 10.810 6.890 ;
        RECT 14.080 6.840 14.460 6.890 ;
        RECT 11.730 0.510 12.020 5.800 ;
        RECT 12.360 0.510 12.530 5.380 ;
        RECT 12.870 0.510 13.160 5.800 ;
        RECT 15.055 0.750 15.355 13.340 ;
        RECT 17.250 8.300 17.540 13.750 ;
        RECT 15.950 7.250 16.330 7.300 ;
        RECT 15.950 6.890 17.280 7.250 ;
        RECT 15.950 6.840 16.330 6.890 ;
        RECT 17.250 0.510 17.540 5.800 ;
        RECT 17.880 0.510 18.050 5.380 ;
        RECT 18.390 0.750 18.690 13.340 ;
        RECT 20.590 8.300 20.880 13.750 ;
        RECT 19.290 7.250 19.670 7.300 ;
        RECT 19.290 6.890 20.620 7.250 ;
        RECT 19.290 6.840 19.670 6.890 ;
        RECT 20.590 0.510 20.880 5.810 ;
        RECT 21.720 0.750 22.020 13.340 ;
        RECT 23.920 8.300 24.210 13.750 ;
        RECT 25.060 8.300 25.350 13.750 ;
        RECT 22.620 7.250 23.000 7.300 ;
        RECT 26.270 7.250 26.650 7.300 ;
        RECT 22.620 6.890 23.950 7.250 ;
        RECT 25.320 6.890 26.650 7.250 ;
        RECT 22.620 6.840 23.000 6.890 ;
        RECT 26.270 6.840 26.650 6.890 ;
        RECT 23.920 0.510 24.210 5.810 ;
        RECT 24.550 0.510 24.720 5.380 ;
        RECT 25.060 0.510 25.350 5.800 ;
        RECT 27.245 0.750 27.545 13.340 ;
        RECT 29.440 8.300 29.730 13.750 ;
        RECT 30.580 8.300 30.870 13.750 ;
        RECT 28.140 7.250 28.520 7.300 ;
        RECT 31.790 7.250 32.170 7.300 ;
        RECT 28.140 6.890 29.470 7.250 ;
        RECT 30.840 6.890 32.170 7.250 ;
        RECT 28.140 6.840 28.520 6.890 ;
        RECT 31.790 6.840 32.170 6.890 ;
        RECT 29.440 0.510 29.730 5.800 ;
        RECT 30.070 0.510 30.240 5.380 ;
        RECT 30.580 0.510 30.870 5.800 ;
        RECT 32.765 0.750 33.065 13.340 ;
        RECT 34.960 8.300 35.250 13.750 ;
        RECT 33.660 7.250 34.040 7.300 ;
        RECT 33.660 6.890 34.990 7.250 ;
        RECT 33.660 6.840 34.040 6.890 ;
        RECT 34.960 0.510 35.250 5.800 ;
        RECT 35.590 0.510 35.760 5.380 ;
        RECT 36.100 0.750 36.400 13.340 ;
        RECT 38.300 8.300 38.590 13.750 ;
        RECT 37.000 7.250 37.380 7.300 ;
        RECT 37.000 6.890 38.330 7.250 ;
        RECT 37.000 6.840 37.380 6.890 ;
        RECT 38.300 0.510 38.590 5.810 ;
        RECT 39.430 0.750 39.730 13.340 ;
        RECT 41.630 8.300 41.920 13.750 ;
        RECT 42.770 8.300 43.060 13.750 ;
        RECT 40.330 7.250 40.710 7.300 ;
        RECT 43.980 7.250 44.360 7.300 ;
        RECT 40.330 6.890 41.660 7.250 ;
        RECT 43.030 6.890 44.360 7.250 ;
        RECT 40.330 6.840 40.710 6.890 ;
        RECT 43.980 6.840 44.360 6.890 ;
        RECT 41.630 0.510 41.920 5.810 ;
        RECT 42.260 0.510 42.430 5.380 ;
        RECT 42.770 0.510 43.060 5.800 ;
        RECT 44.955 0.750 45.255 13.340 ;
        RECT 47.150 8.300 47.440 13.750 ;
        RECT 48.290 8.300 48.580 13.750 ;
        RECT 45.850 7.250 46.230 7.300 ;
        RECT 49.500 7.250 49.880 7.300 ;
        RECT 45.850 6.890 47.180 7.250 ;
        RECT 48.550 6.890 49.880 7.250 ;
        RECT 45.850 6.840 46.230 6.890 ;
        RECT 49.500 6.840 49.880 6.890 ;
        RECT 47.150 0.510 47.440 5.800 ;
        RECT 47.780 0.510 47.950 5.380 ;
        RECT 48.290 0.510 48.580 5.800 ;
        RECT 50.475 0.750 50.775 13.340 ;
        RECT 52.670 8.300 52.960 13.750 ;
        RECT 51.370 7.250 51.750 7.300 ;
        RECT 51.370 6.890 52.700 7.250 ;
        RECT 51.370 6.840 51.750 6.890 ;
        RECT 52.670 0.510 52.960 5.800 ;
        RECT 53.300 0.510 53.470 5.380 ;
        RECT 53.810 0.750 54.110 13.340 ;
        RECT 56.010 8.300 56.300 13.750 ;
        RECT 54.710 7.250 55.090 7.300 ;
        RECT 54.710 6.890 56.040 7.250 ;
        RECT 54.710 6.840 55.090 6.890 ;
        RECT 56.010 0.510 56.300 5.810 ;
        RECT 57.140 0.750 57.440 13.340 ;
        RECT 59.340 8.300 59.630 13.750 ;
        RECT 60.480 8.300 60.770 13.750 ;
        RECT 58.040 7.250 58.420 7.300 ;
        RECT 61.690 7.250 62.070 7.300 ;
        RECT 58.040 6.890 59.370 7.250 ;
        RECT 60.740 6.890 62.070 7.250 ;
        RECT 58.040 6.840 58.420 6.890 ;
        RECT 61.690 6.840 62.070 6.890 ;
        RECT 59.340 0.510 59.630 5.810 ;
        RECT 59.970 0.510 60.140 5.380 ;
        RECT 60.480 0.510 60.770 5.800 ;
        RECT 62.665 0.750 62.965 13.340 ;
        RECT 64.860 8.300 65.150 13.750 ;
        RECT 66.000 8.300 66.290 13.750 ;
        RECT 63.560 7.250 63.940 7.300 ;
        RECT 67.210 7.250 67.590 7.300 ;
        RECT 63.560 6.890 64.890 7.250 ;
        RECT 66.260 6.890 67.590 7.250 ;
        RECT 63.560 6.840 63.940 6.890 ;
        RECT 67.210 6.840 67.590 6.890 ;
        RECT 64.860 0.510 65.150 5.800 ;
        RECT 65.490 0.510 65.660 5.380 ;
        RECT 66.000 0.510 66.290 5.800 ;
        RECT 68.185 0.750 68.485 13.340 ;
        RECT 70.380 8.300 70.670 13.750 ;
        RECT 69.080 7.250 69.460 7.300 ;
        RECT 69.080 6.890 70.410 7.250 ;
        RECT 69.080 6.840 69.460 6.890 ;
        RECT 70.380 0.510 70.670 5.800 ;
        RECT 71.010 0.510 71.180 5.380 ;
        RECT 71.520 0.750 71.820 13.340 ;
        RECT 73.720 8.300 74.010 13.750 ;
        RECT 72.420 7.250 72.800 7.300 ;
        RECT 72.420 6.890 73.750 7.250 ;
        RECT 72.420 6.840 72.800 6.890 ;
        RECT 73.720 0.510 74.010 5.810 ;
        RECT 74.850 0.750 75.150 13.340 ;
        RECT 77.050 8.300 77.340 13.750 ;
        RECT 78.190 8.300 78.480 13.750 ;
        RECT 75.750 7.250 76.130 7.300 ;
        RECT 79.400 7.250 79.780 7.300 ;
        RECT 75.750 6.890 77.080 7.250 ;
        RECT 78.450 6.890 79.780 7.250 ;
        RECT 75.750 6.840 76.130 6.890 ;
        RECT 79.400 6.840 79.780 6.890 ;
        RECT 77.050 0.510 77.340 5.810 ;
        RECT 77.680 0.510 77.850 5.380 ;
        RECT 78.190 0.510 78.480 5.800 ;
        RECT 80.375 0.750 80.675 13.340 ;
        RECT 82.570 8.300 82.860 13.750 ;
        RECT 83.710 8.300 84.000 13.750 ;
        RECT 81.270 7.250 81.650 7.300 ;
        RECT 84.920 7.250 85.300 7.300 ;
        RECT 81.270 6.890 82.600 7.250 ;
        RECT 83.970 6.890 85.300 7.250 ;
        RECT 81.270 6.840 81.650 6.890 ;
        RECT 84.920 6.840 85.300 6.890 ;
        RECT 82.570 0.510 82.860 5.800 ;
        RECT 83.200 0.510 83.370 5.380 ;
        RECT 83.710 0.510 84.000 5.800 ;
        RECT 85.895 0.750 86.195 13.340 ;
        RECT 88.090 8.300 88.380 13.750 ;
        RECT 86.790 7.250 87.170 7.300 ;
        RECT 86.790 6.890 88.120 7.250 ;
        RECT 86.790 6.840 87.170 6.890 ;
        RECT 88.090 0.510 88.380 5.800 ;
        RECT 88.720 0.510 88.890 5.380 ;
        RECT 89.230 0.750 89.530 13.340 ;
        RECT 91.430 8.300 91.720 13.750 ;
        RECT 90.130 7.250 90.510 7.300 ;
        RECT 90.130 6.890 91.460 7.250 ;
        RECT 90.130 6.840 90.510 6.890 ;
        RECT 91.430 0.510 91.720 5.810 ;
        RECT 92.560 0.750 92.860 13.340 ;
        RECT 94.760 8.300 95.050 13.750 ;
        RECT 95.900 8.300 96.190 13.750 ;
        RECT 93.460 7.250 93.840 7.300 ;
        RECT 97.110 7.250 97.490 7.300 ;
        RECT 93.460 6.890 94.790 7.250 ;
        RECT 96.160 6.890 97.490 7.250 ;
        RECT 93.460 6.840 93.840 6.890 ;
        RECT 97.110 6.840 97.490 6.890 ;
        RECT 94.760 0.510 95.050 5.810 ;
        RECT 95.390 0.510 95.560 5.380 ;
        RECT 95.900 0.510 96.190 5.800 ;
        RECT 98.085 0.750 98.385 13.340 ;
        RECT 100.280 8.300 100.570 13.750 ;
        RECT 101.420 8.300 101.710 13.750 ;
        RECT 98.980 7.250 99.360 7.300 ;
        RECT 102.630 7.250 103.010 7.300 ;
        RECT 98.980 6.890 100.310 7.250 ;
        RECT 101.680 6.890 103.010 7.250 ;
        RECT 98.980 6.840 99.360 6.890 ;
        RECT 102.630 6.840 103.010 6.890 ;
        RECT 100.280 0.510 100.570 5.800 ;
        RECT 100.910 0.510 101.080 5.380 ;
        RECT 101.420 0.510 101.710 5.800 ;
        RECT 103.605 0.750 103.905 13.340 ;
        RECT 105.800 8.300 106.090 13.750 ;
        RECT 104.500 7.250 104.880 7.300 ;
        RECT 104.500 6.890 105.830 7.250 ;
        RECT 104.500 6.840 104.880 6.890 ;
        RECT 105.800 0.510 106.090 5.800 ;
        RECT 106.430 0.510 106.600 5.380 ;
        RECT 1.770 0.350 3.170 0.510 ;
        RECT 5.010 0.350 8.860 0.510 ;
        RECT 10.520 0.350 14.370 0.510 ;
        RECT 16.160 0.350 18.050 0.510 ;
        RECT 19.480 0.350 20.880 0.510 ;
        RECT 22.720 0.350 26.570 0.510 ;
        RECT 28.230 0.350 32.080 0.510 ;
        RECT 33.870 0.350 35.760 0.510 ;
        RECT 37.190 0.350 38.590 0.510 ;
        RECT 40.430 0.350 44.280 0.510 ;
        RECT 45.940 0.350 49.790 0.510 ;
        RECT 51.580 0.350 53.470 0.510 ;
        RECT 54.900 0.350 56.300 0.510 ;
        RECT 58.140 0.350 61.990 0.510 ;
        RECT 63.650 0.350 67.500 0.510 ;
        RECT 69.290 0.350 71.180 0.510 ;
        RECT 72.610 0.350 74.010 0.510 ;
        RECT 75.850 0.350 79.700 0.510 ;
        RECT 81.360 0.350 85.210 0.510 ;
        RECT 87.000 0.350 88.890 0.510 ;
        RECT 90.320 0.350 91.720 0.510 ;
        RECT 93.560 0.350 97.410 0.510 ;
        RECT 99.070 0.350 102.920 0.510 ;
        RECT 104.710 0.350 106.600 0.510 ;
        RECT 0.180 0.180 106.600 0.350 ;
        RECT 1.770 0.150 3.170 0.180 ;
        RECT 5.010 0.150 8.860 0.180 ;
        RECT 10.520 0.150 14.370 0.180 ;
        RECT 16.160 0.150 18.050 0.180 ;
        RECT 19.480 0.150 20.880 0.180 ;
        RECT 22.720 0.150 26.570 0.180 ;
        RECT 28.230 0.150 32.080 0.180 ;
        RECT 33.870 0.150 35.760 0.180 ;
        RECT 37.190 0.150 38.590 0.180 ;
        RECT 40.430 0.150 44.280 0.180 ;
        RECT 45.940 0.150 49.790 0.180 ;
        RECT 51.580 0.150 53.470 0.180 ;
        RECT 54.900 0.150 56.300 0.180 ;
        RECT 58.140 0.150 61.990 0.180 ;
        RECT 63.650 0.150 67.500 0.180 ;
        RECT 69.290 0.150 71.180 0.180 ;
        RECT 72.610 0.150 74.010 0.180 ;
        RECT 75.850 0.150 79.700 0.180 ;
        RECT 81.360 0.150 85.210 0.180 ;
        RECT 87.000 0.150 88.890 0.180 ;
        RECT 90.320 0.150 91.720 0.180 ;
        RECT 93.560 0.150 97.410 0.180 ;
        RECT 99.070 0.150 102.920 0.180 ;
        RECT 104.710 0.150 106.600 0.180 ;
      LAYER mcon ;
        RECT 8.720 29.360 9.020 29.660 ;
        RECT 9.210 29.360 9.510 29.660 ;
        RECT 9.700 29.360 10.000 29.660 ;
        RECT 10.190 29.360 10.490 29.660 ;
        RECT 12.400 29.360 12.700 29.660 ;
        RECT 12.890 29.360 13.190 29.660 ;
        RECT 13.380 29.360 13.680 29.660 ;
        RECT 13.870 29.360 14.170 29.660 ;
        RECT 14.360 29.360 14.660 29.660 ;
        RECT 14.850 29.360 15.150 29.660 ;
        RECT 15.340 29.360 15.640 29.660 ;
        RECT 15.830 29.360 16.130 29.660 ;
        RECT 17.910 29.360 18.210 29.660 ;
        RECT 18.400 29.360 18.700 29.660 ;
        RECT 18.890 29.360 19.190 29.660 ;
        RECT 19.380 29.360 19.680 29.660 ;
        RECT 19.870 29.360 20.170 29.660 ;
        RECT 20.360 29.360 20.660 29.660 ;
        RECT 20.850 29.360 21.150 29.660 ;
        RECT 21.340 29.360 21.640 29.660 ;
        RECT 23.600 29.360 23.900 29.660 ;
        RECT 24.090 29.360 24.390 29.660 ;
        RECT 24.580 29.360 24.880 29.660 ;
        RECT 26.430 29.360 26.730 29.660 ;
        RECT 26.920 29.360 27.220 29.660 ;
        RECT 27.410 29.360 27.710 29.660 ;
        RECT 27.900 29.360 28.200 29.660 ;
        RECT 30.110 29.360 30.410 29.660 ;
        RECT 30.600 29.360 30.900 29.660 ;
        RECT 31.090 29.360 31.390 29.660 ;
        RECT 31.580 29.360 31.880 29.660 ;
        RECT 32.070 29.360 32.370 29.660 ;
        RECT 32.560 29.360 32.860 29.660 ;
        RECT 33.050 29.360 33.350 29.660 ;
        RECT 33.540 29.360 33.840 29.660 ;
        RECT 35.620 29.360 35.920 29.660 ;
        RECT 36.110 29.360 36.410 29.660 ;
        RECT 36.600 29.360 36.900 29.660 ;
        RECT 37.090 29.360 37.390 29.660 ;
        RECT 37.580 29.360 37.880 29.660 ;
        RECT 38.070 29.360 38.370 29.660 ;
        RECT 38.560 29.360 38.860 29.660 ;
        RECT 39.050 29.360 39.350 29.660 ;
        RECT 41.310 29.360 41.610 29.660 ;
        RECT 41.800 29.360 42.100 29.660 ;
        RECT 42.290 29.360 42.590 29.660 ;
        RECT 44.140 29.360 44.440 29.660 ;
        RECT 44.630 29.360 44.930 29.660 ;
        RECT 45.120 29.360 45.420 29.660 ;
        RECT 45.610 29.360 45.910 29.660 ;
        RECT 47.820 29.360 48.120 29.660 ;
        RECT 48.310 29.360 48.610 29.660 ;
        RECT 48.800 29.360 49.100 29.660 ;
        RECT 49.290 29.360 49.590 29.660 ;
        RECT 49.780 29.360 50.080 29.660 ;
        RECT 50.270 29.360 50.570 29.660 ;
        RECT 50.760 29.360 51.060 29.660 ;
        RECT 51.250 29.360 51.550 29.660 ;
        RECT 53.330 29.360 53.630 29.660 ;
        RECT 53.820 29.360 54.120 29.660 ;
        RECT 54.310 29.360 54.610 29.660 ;
        RECT 54.800 29.360 55.100 29.660 ;
        RECT 55.290 29.360 55.590 29.660 ;
        RECT 55.780 29.360 56.080 29.660 ;
        RECT 56.270 29.360 56.570 29.660 ;
        RECT 56.760 29.360 57.060 29.660 ;
        RECT 59.020 29.360 59.320 29.660 ;
        RECT 59.510 29.360 59.810 29.660 ;
        RECT 60.000 29.360 60.300 29.660 ;
        RECT 61.850 29.360 62.150 29.660 ;
        RECT 62.340 29.360 62.640 29.660 ;
        RECT 62.830 29.360 63.130 29.660 ;
        RECT 63.320 29.360 63.620 29.660 ;
        RECT 65.530 29.360 65.830 29.660 ;
        RECT 66.020 29.360 66.320 29.660 ;
        RECT 66.510 29.360 66.810 29.660 ;
        RECT 67.000 29.360 67.300 29.660 ;
        RECT 67.490 29.360 67.790 29.660 ;
        RECT 67.980 29.360 68.280 29.660 ;
        RECT 68.470 29.360 68.770 29.660 ;
        RECT 68.960 29.360 69.260 29.660 ;
        RECT 71.040 29.360 71.340 29.660 ;
        RECT 71.530 29.360 71.830 29.660 ;
        RECT 72.020 29.360 72.320 29.660 ;
        RECT 72.510 29.360 72.810 29.660 ;
        RECT 73.000 29.360 73.300 29.660 ;
        RECT 73.490 29.360 73.790 29.660 ;
        RECT 73.980 29.360 74.280 29.660 ;
        RECT 74.470 29.360 74.770 29.660 ;
        RECT 76.730 29.360 77.030 29.660 ;
        RECT 77.220 29.360 77.520 29.660 ;
        RECT 77.710 29.360 78.010 29.660 ;
        RECT 79.560 29.360 79.860 29.660 ;
        RECT 80.050 29.360 80.350 29.660 ;
        RECT 80.540 29.360 80.840 29.660 ;
        RECT 81.030 29.360 81.330 29.660 ;
        RECT 83.240 29.360 83.540 29.660 ;
        RECT 83.730 29.360 84.030 29.660 ;
        RECT 84.220 29.360 84.520 29.660 ;
        RECT 84.710 29.360 85.010 29.660 ;
        RECT 85.200 29.360 85.500 29.660 ;
        RECT 85.690 29.360 85.990 29.660 ;
        RECT 86.180 29.360 86.480 29.660 ;
        RECT 86.670 29.360 86.970 29.660 ;
        RECT 88.750 29.360 89.050 29.660 ;
        RECT 89.240 29.360 89.540 29.660 ;
        RECT 89.730 29.360 90.030 29.660 ;
        RECT 90.220 29.360 90.520 29.660 ;
        RECT 90.710 29.360 91.010 29.660 ;
        RECT 91.200 29.360 91.500 29.660 ;
        RECT 91.690 29.360 91.990 29.660 ;
        RECT 92.180 29.360 92.480 29.660 ;
        RECT 94.440 29.360 94.740 29.660 ;
        RECT 94.930 29.360 95.230 29.660 ;
        RECT 95.420 29.360 95.720 29.660 ;
        RECT -0.665 25.435 -0.495 25.605 ;
        RECT -0.205 25.435 -0.035 25.605 ;
        RECT 0.255 25.435 0.425 25.605 ;
        RECT 0.715 25.435 0.885 25.605 ;
        RECT 1.175 25.435 1.345 25.605 ;
        RECT 3.330 25.435 3.500 25.605 ;
        RECT 3.790 25.435 3.960 25.605 ;
        RECT 4.250 25.435 4.420 25.605 ;
        RECT 2.240 24.040 2.480 24.280 ;
        RECT 11.355 23.980 11.655 24.280 ;
        RECT -0.665 22.715 -0.495 22.885 ;
        RECT -0.205 22.715 -0.035 22.885 ;
        RECT 0.255 22.715 0.425 22.885 ;
        RECT 0.715 22.715 0.885 22.885 ;
        RECT 1.175 22.715 1.345 22.885 ;
        RECT 3.330 22.715 3.500 22.885 ;
        RECT 3.790 22.715 3.960 22.885 ;
        RECT 4.250 22.715 4.420 22.885 ;
        RECT 9.430 22.620 9.730 22.920 ;
        RECT 9.920 22.620 10.220 22.920 ;
        RECT 10.410 22.620 10.710 22.920 ;
        RECT 12.300 22.620 12.600 22.920 ;
        RECT 12.790 22.620 13.090 22.920 ;
        RECT 13.280 22.620 13.580 22.920 ;
        RECT 14.950 22.620 15.250 22.920 ;
        RECT 15.440 22.620 15.740 22.920 ;
        RECT 15.930 22.620 16.230 22.920 ;
        RECT 17.820 22.620 18.120 22.920 ;
        RECT 18.310 22.620 18.610 22.920 ;
        RECT 18.800 22.620 19.100 22.920 ;
        RECT 20.470 22.620 20.770 22.920 ;
        RECT 20.960 22.620 21.260 22.920 ;
        RECT 21.450 22.620 21.750 22.920 ;
        RECT 16.875 21.260 17.175 21.560 ;
        RECT 25.730 23.980 26.030 24.280 ;
        RECT 23.800 22.620 24.100 22.920 ;
        RECT 24.290 22.620 24.590 22.920 ;
        RECT 24.780 22.620 25.080 22.920 ;
        RECT 22.400 21.260 22.700 21.560 ;
        RECT 29.065 23.980 29.365 24.280 ;
        RECT 27.140 22.620 27.440 22.920 ;
        RECT 27.630 22.620 27.930 22.920 ;
        RECT 28.120 22.620 28.420 22.920 ;
        RECT 30.010 22.620 30.310 22.920 ;
        RECT 30.500 22.620 30.800 22.920 ;
        RECT 30.990 22.620 31.290 22.920 ;
        RECT 32.660 22.620 32.960 22.920 ;
        RECT 33.150 22.620 33.450 22.920 ;
        RECT 33.640 22.620 33.940 22.920 ;
        RECT 35.530 22.620 35.830 22.920 ;
        RECT 36.020 22.620 36.320 22.920 ;
        RECT 36.510 22.620 36.810 22.920 ;
        RECT 38.180 22.620 38.480 22.920 ;
        RECT 38.670 22.620 38.970 22.920 ;
        RECT 39.160 22.620 39.460 22.920 ;
        RECT 34.585 21.260 34.885 21.560 ;
        RECT 43.440 23.980 43.740 24.280 ;
        RECT 41.510 22.620 41.810 22.920 ;
        RECT 42.000 22.620 42.300 22.920 ;
        RECT 42.490 22.620 42.790 22.920 ;
        RECT 40.110 21.260 40.410 21.560 ;
        RECT 46.775 23.980 47.075 24.280 ;
        RECT 44.850 22.620 45.150 22.920 ;
        RECT 45.340 22.620 45.640 22.920 ;
        RECT 45.830 22.620 46.130 22.920 ;
        RECT 47.720 22.620 48.020 22.920 ;
        RECT 48.210 22.620 48.510 22.920 ;
        RECT 48.700 22.620 49.000 22.920 ;
        RECT 50.370 22.620 50.670 22.920 ;
        RECT 50.860 22.620 51.160 22.920 ;
        RECT 51.350 22.620 51.650 22.920 ;
        RECT 53.240 22.620 53.540 22.920 ;
        RECT 53.730 22.620 54.030 22.920 ;
        RECT 54.220 22.620 54.520 22.920 ;
        RECT 55.890 22.620 56.190 22.920 ;
        RECT 56.380 22.620 56.680 22.920 ;
        RECT 56.870 22.620 57.170 22.920 ;
        RECT 52.295 21.260 52.595 21.560 ;
        RECT 61.150 23.980 61.450 24.280 ;
        RECT 59.220 22.620 59.520 22.920 ;
        RECT 59.710 22.620 60.010 22.920 ;
        RECT 60.200 22.620 60.500 22.920 ;
        RECT 57.820 21.260 58.120 21.560 ;
        RECT 64.485 23.980 64.785 24.280 ;
        RECT 62.560 22.620 62.860 22.920 ;
        RECT 63.050 22.620 63.350 22.920 ;
        RECT 63.540 22.620 63.840 22.920 ;
        RECT 65.430 22.620 65.730 22.920 ;
        RECT 65.920 22.620 66.220 22.920 ;
        RECT 66.410 22.620 66.710 22.920 ;
        RECT 68.080 22.620 68.380 22.920 ;
        RECT 68.570 22.620 68.870 22.920 ;
        RECT 69.060 22.620 69.360 22.920 ;
        RECT 70.950 22.620 71.250 22.920 ;
        RECT 71.440 22.620 71.740 22.920 ;
        RECT 71.930 22.620 72.230 22.920 ;
        RECT 73.600 22.620 73.900 22.920 ;
        RECT 74.090 22.620 74.390 22.920 ;
        RECT 74.580 22.620 74.880 22.920 ;
        RECT 70.005 21.260 70.305 21.560 ;
        RECT 78.860 23.980 79.160 24.280 ;
        RECT 76.930 22.620 77.230 22.920 ;
        RECT 77.420 22.620 77.720 22.920 ;
        RECT 77.910 22.620 78.210 22.920 ;
        RECT 75.530 21.260 75.830 21.560 ;
        RECT 82.195 23.980 82.495 24.280 ;
        RECT 80.270 22.620 80.570 22.920 ;
        RECT 80.760 22.620 81.060 22.920 ;
        RECT 81.250 22.620 81.550 22.920 ;
        RECT 83.140 22.620 83.440 22.920 ;
        RECT 83.630 22.620 83.930 22.920 ;
        RECT 84.120 22.620 84.420 22.920 ;
        RECT 85.790 22.620 86.090 22.920 ;
        RECT 86.280 22.620 86.580 22.920 ;
        RECT 86.770 22.620 87.070 22.920 ;
        RECT 88.660 22.620 88.960 22.920 ;
        RECT 89.150 22.620 89.450 22.920 ;
        RECT 89.640 22.620 89.940 22.920 ;
        RECT 91.310 22.620 91.610 22.920 ;
        RECT 91.800 22.620 92.100 22.920 ;
        RECT 92.290 22.620 92.590 22.920 ;
        RECT 87.715 21.260 88.015 21.560 ;
        RECT 96.570 23.980 96.870 24.280 ;
        RECT 101.100 24.050 101.400 24.350 ;
        RECT 101.600 24.050 101.900 24.350 ;
        RECT 102.100 24.050 102.400 24.350 ;
        RECT 102.600 24.050 102.900 24.350 ;
        RECT 94.640 22.620 94.940 22.920 ;
        RECT 95.130 22.620 95.430 22.920 ;
        RECT 95.620 22.620 95.920 22.920 ;
        RECT 93.240 21.260 93.540 21.560 ;
        RECT 102.090 19.120 102.390 19.420 ;
        RECT 102.610 19.120 102.910 19.420 ;
        RECT 102.090 18.600 102.390 18.900 ;
        RECT 102.610 18.600 102.910 18.900 ;
        RECT 107.605 19.100 107.905 19.400 ;
        RECT 108.095 19.100 108.395 19.400 ;
        RECT 107.605 18.600 107.905 18.900 ;
        RECT 108.095 18.600 108.395 18.900 ;
        RECT 8.720 15.760 9.020 16.060 ;
        RECT 9.210 15.760 9.510 16.060 ;
        RECT 9.700 15.760 10.000 16.060 ;
        RECT 10.190 15.760 10.490 16.060 ;
        RECT 12.400 15.760 12.700 16.060 ;
        RECT 12.890 15.760 13.190 16.060 ;
        RECT 13.380 15.760 13.680 16.060 ;
        RECT 13.870 15.760 14.170 16.060 ;
        RECT 14.360 15.760 14.660 16.060 ;
        RECT 14.850 15.760 15.150 16.060 ;
        RECT 15.340 15.760 15.640 16.060 ;
        RECT 15.830 15.760 16.130 16.060 ;
        RECT 17.910 15.760 18.210 16.060 ;
        RECT 18.400 15.760 18.700 16.060 ;
        RECT 18.890 15.760 19.190 16.060 ;
        RECT 19.380 15.760 19.680 16.060 ;
        RECT 19.870 15.760 20.170 16.060 ;
        RECT 20.360 15.760 20.660 16.060 ;
        RECT 20.850 15.760 21.150 16.060 ;
        RECT 21.340 15.760 21.640 16.060 ;
        RECT 23.600 15.760 23.900 16.060 ;
        RECT 24.090 15.760 24.390 16.060 ;
        RECT 24.580 15.760 24.880 16.060 ;
        RECT 26.430 15.760 26.730 16.060 ;
        RECT 26.920 15.760 27.220 16.060 ;
        RECT 27.410 15.760 27.710 16.060 ;
        RECT 27.900 15.760 28.200 16.060 ;
        RECT 30.110 15.760 30.410 16.060 ;
        RECT 30.600 15.760 30.900 16.060 ;
        RECT 31.090 15.760 31.390 16.060 ;
        RECT 31.580 15.760 31.880 16.060 ;
        RECT 32.070 15.760 32.370 16.060 ;
        RECT 32.560 15.760 32.860 16.060 ;
        RECT 33.050 15.760 33.350 16.060 ;
        RECT 33.540 15.760 33.840 16.060 ;
        RECT 35.620 15.760 35.920 16.060 ;
        RECT 36.110 15.760 36.410 16.060 ;
        RECT 36.600 15.760 36.900 16.060 ;
        RECT 37.090 15.760 37.390 16.060 ;
        RECT 37.580 15.760 37.880 16.060 ;
        RECT 38.070 15.760 38.370 16.060 ;
        RECT 38.560 15.760 38.860 16.060 ;
        RECT 39.050 15.760 39.350 16.060 ;
        RECT 41.310 15.760 41.610 16.060 ;
        RECT 41.800 15.760 42.100 16.060 ;
        RECT 42.290 15.760 42.590 16.060 ;
        RECT 44.140 15.760 44.440 16.060 ;
        RECT 44.630 15.760 44.930 16.060 ;
        RECT 45.120 15.760 45.420 16.060 ;
        RECT 45.610 15.760 45.910 16.060 ;
        RECT 47.820 15.760 48.120 16.060 ;
        RECT 48.310 15.760 48.610 16.060 ;
        RECT 48.800 15.760 49.100 16.060 ;
        RECT 49.290 15.760 49.590 16.060 ;
        RECT 49.780 15.760 50.080 16.060 ;
        RECT 50.270 15.760 50.570 16.060 ;
        RECT 50.760 15.760 51.060 16.060 ;
        RECT 51.250 15.760 51.550 16.060 ;
        RECT 53.330 15.760 53.630 16.060 ;
        RECT 53.820 15.760 54.120 16.060 ;
        RECT 54.310 15.760 54.610 16.060 ;
        RECT 54.800 15.760 55.100 16.060 ;
        RECT 55.290 15.760 55.590 16.060 ;
        RECT 55.780 15.760 56.080 16.060 ;
        RECT 56.270 15.760 56.570 16.060 ;
        RECT 56.760 15.760 57.060 16.060 ;
        RECT 59.020 15.760 59.320 16.060 ;
        RECT 59.510 15.760 59.810 16.060 ;
        RECT 60.000 15.760 60.300 16.060 ;
        RECT 61.850 15.760 62.150 16.060 ;
        RECT 62.340 15.760 62.640 16.060 ;
        RECT 62.830 15.760 63.130 16.060 ;
        RECT 63.320 15.760 63.620 16.060 ;
        RECT 65.530 15.760 65.830 16.060 ;
        RECT 66.020 15.760 66.320 16.060 ;
        RECT 66.510 15.760 66.810 16.060 ;
        RECT 67.000 15.760 67.300 16.060 ;
        RECT 67.490 15.760 67.790 16.060 ;
        RECT 67.980 15.760 68.280 16.060 ;
        RECT 68.470 15.760 68.770 16.060 ;
        RECT 68.960 15.760 69.260 16.060 ;
        RECT 71.040 15.760 71.340 16.060 ;
        RECT 71.530 15.760 71.830 16.060 ;
        RECT 72.020 15.760 72.320 16.060 ;
        RECT 72.510 15.760 72.810 16.060 ;
        RECT 73.000 15.760 73.300 16.060 ;
        RECT 73.490 15.760 73.790 16.060 ;
        RECT 73.980 15.760 74.280 16.060 ;
        RECT 74.470 15.760 74.770 16.060 ;
        RECT 76.730 15.760 77.030 16.060 ;
        RECT 77.220 15.760 77.520 16.060 ;
        RECT 77.710 15.760 78.010 16.060 ;
        RECT 79.560 15.760 79.860 16.060 ;
        RECT 80.050 15.760 80.350 16.060 ;
        RECT 80.540 15.760 80.840 16.060 ;
        RECT 81.030 15.760 81.330 16.060 ;
        RECT 83.240 15.760 83.540 16.060 ;
        RECT 83.730 15.760 84.030 16.060 ;
        RECT 84.220 15.760 84.520 16.060 ;
        RECT 84.710 15.760 85.010 16.060 ;
        RECT 85.200 15.760 85.500 16.060 ;
        RECT 85.690 15.760 85.990 16.060 ;
        RECT 86.180 15.760 86.480 16.060 ;
        RECT 86.670 15.760 86.970 16.060 ;
        RECT 88.750 15.760 89.050 16.060 ;
        RECT 89.240 15.760 89.540 16.060 ;
        RECT 89.730 15.760 90.030 16.060 ;
        RECT 90.220 15.760 90.520 16.060 ;
        RECT 90.710 15.760 91.010 16.060 ;
        RECT 91.200 15.760 91.500 16.060 ;
        RECT 91.690 15.760 91.990 16.060 ;
        RECT 92.180 15.760 92.480 16.060 ;
        RECT 94.440 15.760 94.740 16.060 ;
        RECT 94.930 15.760 95.230 16.060 ;
        RECT 95.420 15.760 95.720 16.060 ;
        RECT 1.830 13.780 2.130 14.080 ;
        RECT 2.320 13.780 2.620 14.080 ;
        RECT 2.810 13.780 3.110 14.080 ;
        RECT 5.070 13.780 5.370 14.080 ;
        RECT 5.560 13.780 5.860 14.080 ;
        RECT 6.050 13.780 6.350 14.080 ;
        RECT 6.540 13.780 6.840 14.080 ;
        RECT 7.030 13.780 7.330 14.080 ;
        RECT 7.520 13.780 7.820 14.080 ;
        RECT 8.010 13.780 8.310 14.080 ;
        RECT 8.500 13.780 8.800 14.080 ;
        RECT 10.580 13.780 10.880 14.080 ;
        RECT 11.070 13.780 11.370 14.080 ;
        RECT 11.560 13.780 11.860 14.080 ;
        RECT 12.050 13.780 12.350 14.080 ;
        RECT 12.540 13.780 12.840 14.080 ;
        RECT 13.030 13.780 13.330 14.080 ;
        RECT 13.520 13.780 13.820 14.080 ;
        RECT 14.010 13.780 14.310 14.080 ;
        RECT 16.220 13.780 16.520 14.080 ;
        RECT 16.710 13.780 17.010 14.080 ;
        RECT 17.200 13.780 17.500 14.080 ;
        RECT 17.690 13.780 17.990 14.080 ;
        RECT 19.540 13.780 19.840 14.080 ;
        RECT 20.030 13.780 20.330 14.080 ;
        RECT 20.520 13.780 20.820 14.080 ;
        RECT 22.780 13.780 23.080 14.080 ;
        RECT 23.270 13.780 23.570 14.080 ;
        RECT 23.760 13.780 24.060 14.080 ;
        RECT 24.250 13.780 24.550 14.080 ;
        RECT 24.740 13.780 25.040 14.080 ;
        RECT 25.230 13.780 25.530 14.080 ;
        RECT 25.720 13.780 26.020 14.080 ;
        RECT 26.210 13.780 26.510 14.080 ;
        RECT 28.290 13.780 28.590 14.080 ;
        RECT 28.780 13.780 29.080 14.080 ;
        RECT 29.270 13.780 29.570 14.080 ;
        RECT 29.760 13.780 30.060 14.080 ;
        RECT 30.250 13.780 30.550 14.080 ;
        RECT 30.740 13.780 31.040 14.080 ;
        RECT 31.230 13.780 31.530 14.080 ;
        RECT 31.720 13.780 32.020 14.080 ;
        RECT 33.930 13.780 34.230 14.080 ;
        RECT 34.420 13.780 34.720 14.080 ;
        RECT 34.910 13.780 35.210 14.080 ;
        RECT 35.400 13.780 35.700 14.080 ;
        RECT 37.250 13.780 37.550 14.080 ;
        RECT 37.740 13.780 38.040 14.080 ;
        RECT 38.230 13.780 38.530 14.080 ;
        RECT 40.490 13.780 40.790 14.080 ;
        RECT 40.980 13.780 41.280 14.080 ;
        RECT 41.470 13.780 41.770 14.080 ;
        RECT 41.960 13.780 42.260 14.080 ;
        RECT 42.450 13.780 42.750 14.080 ;
        RECT 42.940 13.780 43.240 14.080 ;
        RECT 43.430 13.780 43.730 14.080 ;
        RECT 43.920 13.780 44.220 14.080 ;
        RECT 46.000 13.780 46.300 14.080 ;
        RECT 46.490 13.780 46.790 14.080 ;
        RECT 46.980 13.780 47.280 14.080 ;
        RECT 47.470 13.780 47.770 14.080 ;
        RECT 47.960 13.780 48.260 14.080 ;
        RECT 48.450 13.780 48.750 14.080 ;
        RECT 48.940 13.780 49.240 14.080 ;
        RECT 49.430 13.780 49.730 14.080 ;
        RECT 51.640 13.780 51.940 14.080 ;
        RECT 52.130 13.780 52.430 14.080 ;
        RECT 52.620 13.780 52.920 14.080 ;
        RECT 53.110 13.780 53.410 14.080 ;
        RECT 54.960 13.780 55.260 14.080 ;
        RECT 55.450 13.780 55.750 14.080 ;
        RECT 55.940 13.780 56.240 14.080 ;
        RECT 58.200 13.780 58.500 14.080 ;
        RECT 58.690 13.780 58.990 14.080 ;
        RECT 59.180 13.780 59.480 14.080 ;
        RECT 59.670 13.780 59.970 14.080 ;
        RECT 60.160 13.780 60.460 14.080 ;
        RECT 60.650 13.780 60.950 14.080 ;
        RECT 61.140 13.780 61.440 14.080 ;
        RECT 61.630 13.780 61.930 14.080 ;
        RECT 63.710 13.780 64.010 14.080 ;
        RECT 64.200 13.780 64.500 14.080 ;
        RECT 64.690 13.780 64.990 14.080 ;
        RECT 65.180 13.780 65.480 14.080 ;
        RECT 65.670 13.780 65.970 14.080 ;
        RECT 66.160 13.780 66.460 14.080 ;
        RECT 66.650 13.780 66.950 14.080 ;
        RECT 67.140 13.780 67.440 14.080 ;
        RECT 69.350 13.780 69.650 14.080 ;
        RECT 69.840 13.780 70.140 14.080 ;
        RECT 70.330 13.780 70.630 14.080 ;
        RECT 70.820 13.780 71.120 14.080 ;
        RECT 72.670 13.780 72.970 14.080 ;
        RECT 73.160 13.780 73.460 14.080 ;
        RECT 73.650 13.780 73.950 14.080 ;
        RECT 75.910 13.780 76.210 14.080 ;
        RECT 76.400 13.780 76.700 14.080 ;
        RECT 76.890 13.780 77.190 14.080 ;
        RECT 77.380 13.780 77.680 14.080 ;
        RECT 77.870 13.780 78.170 14.080 ;
        RECT 78.360 13.780 78.660 14.080 ;
        RECT 78.850 13.780 79.150 14.080 ;
        RECT 79.340 13.780 79.640 14.080 ;
        RECT 81.420 13.780 81.720 14.080 ;
        RECT 81.910 13.780 82.210 14.080 ;
        RECT 82.400 13.780 82.700 14.080 ;
        RECT 82.890 13.780 83.190 14.080 ;
        RECT 83.380 13.780 83.680 14.080 ;
        RECT 83.870 13.780 84.170 14.080 ;
        RECT 84.360 13.780 84.660 14.080 ;
        RECT 84.850 13.780 85.150 14.080 ;
        RECT 87.060 13.780 87.360 14.080 ;
        RECT 87.550 13.780 87.850 14.080 ;
        RECT 88.040 13.780 88.340 14.080 ;
        RECT 88.530 13.780 88.830 14.080 ;
        RECT 90.380 13.780 90.680 14.080 ;
        RECT 90.870 13.780 91.170 14.080 ;
        RECT 91.360 13.780 91.660 14.080 ;
        RECT 93.620 13.780 93.920 14.080 ;
        RECT 94.110 13.780 94.410 14.080 ;
        RECT 94.600 13.780 94.900 14.080 ;
        RECT 95.090 13.780 95.390 14.080 ;
        RECT 95.580 13.780 95.880 14.080 ;
        RECT 96.070 13.780 96.370 14.080 ;
        RECT 96.560 13.780 96.860 14.080 ;
        RECT 97.050 13.780 97.350 14.080 ;
        RECT 99.130 13.780 99.430 14.080 ;
        RECT 99.620 13.780 99.920 14.080 ;
        RECT 100.110 13.780 100.410 14.080 ;
        RECT 100.600 13.780 100.900 14.080 ;
        RECT 101.090 13.780 101.390 14.080 ;
        RECT 101.580 13.780 101.880 14.080 ;
        RECT 102.070 13.780 102.370 14.080 ;
        RECT 102.560 13.780 102.860 14.080 ;
        RECT 104.770 13.780 105.070 14.080 ;
        RECT 105.260 13.780 105.560 14.080 ;
        RECT 105.750 13.780 106.050 14.080 ;
        RECT 106.240 13.780 106.540 14.080 ;
        RECT 4.010 8.280 4.310 8.580 ;
        RECT 1.630 6.920 1.930 7.220 ;
        RECT 2.120 6.920 2.420 7.220 ;
        RECT 2.610 6.920 2.910 7.220 ;
        RECT 0.680 5.560 0.980 5.860 ;
        RECT 9.535 8.280 9.835 8.580 ;
        RECT 4.960 6.920 5.260 7.220 ;
        RECT 5.450 6.920 5.750 7.220 ;
        RECT 5.940 6.920 6.240 7.220 ;
        RECT 7.610 6.920 7.910 7.220 ;
        RECT 8.100 6.920 8.400 7.220 ;
        RECT 8.590 6.920 8.890 7.220 ;
        RECT 10.480 6.920 10.780 7.220 ;
        RECT 10.970 6.920 11.270 7.220 ;
        RECT 11.460 6.920 11.760 7.220 ;
        RECT 13.130 6.920 13.430 7.220 ;
        RECT 13.620 6.920 13.920 7.220 ;
        RECT 14.110 6.920 14.410 7.220 ;
        RECT 16.000 6.920 16.300 7.220 ;
        RECT 16.490 6.920 16.790 7.220 ;
        RECT 16.980 6.920 17.280 7.220 ;
        RECT 15.055 5.560 15.355 5.860 ;
        RECT 21.720 8.280 22.020 8.580 ;
        RECT 19.340 6.920 19.640 7.220 ;
        RECT 19.830 6.920 20.130 7.220 ;
        RECT 20.320 6.920 20.620 7.220 ;
        RECT 18.390 5.560 18.690 5.860 ;
        RECT 27.245 8.280 27.545 8.580 ;
        RECT 22.670 6.920 22.970 7.220 ;
        RECT 23.160 6.920 23.460 7.220 ;
        RECT 23.650 6.920 23.950 7.220 ;
        RECT 25.320 6.920 25.620 7.220 ;
        RECT 25.810 6.920 26.110 7.220 ;
        RECT 26.300 6.920 26.600 7.220 ;
        RECT 28.190 6.920 28.490 7.220 ;
        RECT 28.680 6.920 28.980 7.220 ;
        RECT 29.170 6.920 29.470 7.220 ;
        RECT 30.840 6.920 31.140 7.220 ;
        RECT 31.330 6.920 31.630 7.220 ;
        RECT 31.820 6.920 32.120 7.220 ;
        RECT 33.710 6.920 34.010 7.220 ;
        RECT 34.200 6.920 34.500 7.220 ;
        RECT 34.690 6.920 34.990 7.220 ;
        RECT 32.765 5.560 33.065 5.860 ;
        RECT 39.430 8.280 39.730 8.580 ;
        RECT 37.050 6.920 37.350 7.220 ;
        RECT 37.540 6.920 37.840 7.220 ;
        RECT 38.030 6.920 38.330 7.220 ;
        RECT 36.100 5.560 36.400 5.860 ;
        RECT 44.955 8.280 45.255 8.580 ;
        RECT 40.380 6.920 40.680 7.220 ;
        RECT 40.870 6.920 41.170 7.220 ;
        RECT 41.360 6.920 41.660 7.220 ;
        RECT 43.030 6.920 43.330 7.220 ;
        RECT 43.520 6.920 43.820 7.220 ;
        RECT 44.010 6.920 44.310 7.220 ;
        RECT 45.900 6.920 46.200 7.220 ;
        RECT 46.390 6.920 46.690 7.220 ;
        RECT 46.880 6.920 47.180 7.220 ;
        RECT 48.550 6.920 48.850 7.220 ;
        RECT 49.040 6.920 49.340 7.220 ;
        RECT 49.530 6.920 49.830 7.220 ;
        RECT 51.420 6.920 51.720 7.220 ;
        RECT 51.910 6.920 52.210 7.220 ;
        RECT 52.400 6.920 52.700 7.220 ;
        RECT 50.475 5.560 50.775 5.860 ;
        RECT 57.140 8.280 57.440 8.580 ;
        RECT 54.760 6.920 55.060 7.220 ;
        RECT 55.250 6.920 55.550 7.220 ;
        RECT 55.740 6.920 56.040 7.220 ;
        RECT 53.810 5.560 54.110 5.860 ;
        RECT 62.665 8.280 62.965 8.580 ;
        RECT 58.090 6.920 58.390 7.220 ;
        RECT 58.580 6.920 58.880 7.220 ;
        RECT 59.070 6.920 59.370 7.220 ;
        RECT 60.740 6.920 61.040 7.220 ;
        RECT 61.230 6.920 61.530 7.220 ;
        RECT 61.720 6.920 62.020 7.220 ;
        RECT 63.610 6.920 63.910 7.220 ;
        RECT 64.100 6.920 64.400 7.220 ;
        RECT 64.590 6.920 64.890 7.220 ;
        RECT 66.260 6.920 66.560 7.220 ;
        RECT 66.750 6.920 67.050 7.220 ;
        RECT 67.240 6.920 67.540 7.220 ;
        RECT 69.130 6.920 69.430 7.220 ;
        RECT 69.620 6.920 69.920 7.220 ;
        RECT 70.110 6.920 70.410 7.220 ;
        RECT 68.185 5.560 68.485 5.860 ;
        RECT 74.850 8.280 75.150 8.580 ;
        RECT 72.470 6.920 72.770 7.220 ;
        RECT 72.960 6.920 73.260 7.220 ;
        RECT 73.450 6.920 73.750 7.220 ;
        RECT 71.520 5.560 71.820 5.860 ;
        RECT 80.375 8.280 80.675 8.580 ;
        RECT 75.800 6.920 76.100 7.220 ;
        RECT 76.290 6.920 76.590 7.220 ;
        RECT 76.780 6.920 77.080 7.220 ;
        RECT 78.450 6.920 78.750 7.220 ;
        RECT 78.940 6.920 79.240 7.220 ;
        RECT 79.430 6.920 79.730 7.220 ;
        RECT 81.320 6.920 81.620 7.220 ;
        RECT 81.810 6.920 82.110 7.220 ;
        RECT 82.300 6.920 82.600 7.220 ;
        RECT 83.970 6.920 84.270 7.220 ;
        RECT 84.460 6.920 84.760 7.220 ;
        RECT 84.950 6.920 85.250 7.220 ;
        RECT 86.840 6.920 87.140 7.220 ;
        RECT 87.330 6.920 87.630 7.220 ;
        RECT 87.820 6.920 88.120 7.220 ;
        RECT 85.895 5.560 86.195 5.860 ;
        RECT 92.560 8.280 92.860 8.580 ;
        RECT 90.180 6.920 90.480 7.220 ;
        RECT 90.670 6.920 90.970 7.220 ;
        RECT 91.160 6.920 91.460 7.220 ;
        RECT 89.230 5.560 89.530 5.860 ;
        RECT 98.085 8.280 98.385 8.580 ;
        RECT 93.510 6.920 93.810 7.220 ;
        RECT 94.000 6.920 94.300 7.220 ;
        RECT 94.490 6.920 94.790 7.220 ;
        RECT 96.160 6.920 96.460 7.220 ;
        RECT 96.650 6.920 96.950 7.220 ;
        RECT 97.140 6.920 97.440 7.220 ;
        RECT 99.030 6.920 99.330 7.220 ;
        RECT 99.520 6.920 99.820 7.220 ;
        RECT 100.010 6.920 100.310 7.220 ;
        RECT 101.680 6.920 101.980 7.220 ;
        RECT 102.170 6.920 102.470 7.220 ;
        RECT 102.660 6.920 102.960 7.220 ;
        RECT 104.550 6.920 104.850 7.220 ;
        RECT 105.040 6.920 105.340 7.220 ;
        RECT 105.530 6.920 105.830 7.220 ;
        RECT 103.605 5.560 103.905 5.860 ;
        RECT 1.830 0.180 2.130 0.480 ;
        RECT 2.320 0.180 2.620 0.480 ;
        RECT 2.810 0.180 3.110 0.480 ;
        RECT 5.070 0.180 5.370 0.480 ;
        RECT 5.560 0.180 5.860 0.480 ;
        RECT 6.050 0.180 6.350 0.480 ;
        RECT 6.540 0.180 6.840 0.480 ;
        RECT 7.030 0.180 7.330 0.480 ;
        RECT 7.520 0.180 7.820 0.480 ;
        RECT 8.010 0.180 8.310 0.480 ;
        RECT 8.500 0.180 8.800 0.480 ;
        RECT 10.580 0.180 10.880 0.480 ;
        RECT 11.070 0.180 11.370 0.480 ;
        RECT 11.560 0.180 11.860 0.480 ;
        RECT 12.050 0.180 12.350 0.480 ;
        RECT 12.540 0.180 12.840 0.480 ;
        RECT 13.030 0.180 13.330 0.480 ;
        RECT 13.520 0.180 13.820 0.480 ;
        RECT 14.010 0.180 14.310 0.480 ;
        RECT 16.220 0.180 16.520 0.480 ;
        RECT 16.710 0.180 17.010 0.480 ;
        RECT 17.200 0.180 17.500 0.480 ;
        RECT 17.690 0.180 17.990 0.480 ;
        RECT 19.540 0.180 19.840 0.480 ;
        RECT 20.030 0.180 20.330 0.480 ;
        RECT 20.520 0.180 20.820 0.480 ;
        RECT 22.780 0.180 23.080 0.480 ;
        RECT 23.270 0.180 23.570 0.480 ;
        RECT 23.760 0.180 24.060 0.480 ;
        RECT 24.250 0.180 24.550 0.480 ;
        RECT 24.740 0.180 25.040 0.480 ;
        RECT 25.230 0.180 25.530 0.480 ;
        RECT 25.720 0.180 26.020 0.480 ;
        RECT 26.210 0.180 26.510 0.480 ;
        RECT 28.290 0.180 28.590 0.480 ;
        RECT 28.780 0.180 29.080 0.480 ;
        RECT 29.270 0.180 29.570 0.480 ;
        RECT 29.760 0.180 30.060 0.480 ;
        RECT 30.250 0.180 30.550 0.480 ;
        RECT 30.740 0.180 31.040 0.480 ;
        RECT 31.230 0.180 31.530 0.480 ;
        RECT 31.720 0.180 32.020 0.480 ;
        RECT 33.930 0.180 34.230 0.480 ;
        RECT 34.420 0.180 34.720 0.480 ;
        RECT 34.910 0.180 35.210 0.480 ;
        RECT 35.400 0.180 35.700 0.480 ;
        RECT 37.250 0.180 37.550 0.480 ;
        RECT 37.740 0.180 38.040 0.480 ;
        RECT 38.230 0.180 38.530 0.480 ;
        RECT 40.490 0.180 40.790 0.480 ;
        RECT 40.980 0.180 41.280 0.480 ;
        RECT 41.470 0.180 41.770 0.480 ;
        RECT 41.960 0.180 42.260 0.480 ;
        RECT 42.450 0.180 42.750 0.480 ;
        RECT 42.940 0.180 43.240 0.480 ;
        RECT 43.430 0.180 43.730 0.480 ;
        RECT 43.920 0.180 44.220 0.480 ;
        RECT 46.000 0.180 46.300 0.480 ;
        RECT 46.490 0.180 46.790 0.480 ;
        RECT 46.980 0.180 47.280 0.480 ;
        RECT 47.470 0.180 47.770 0.480 ;
        RECT 47.960 0.180 48.260 0.480 ;
        RECT 48.450 0.180 48.750 0.480 ;
        RECT 48.940 0.180 49.240 0.480 ;
        RECT 49.430 0.180 49.730 0.480 ;
        RECT 51.640 0.180 51.940 0.480 ;
        RECT 52.130 0.180 52.430 0.480 ;
        RECT 52.620 0.180 52.920 0.480 ;
        RECT 53.110 0.180 53.410 0.480 ;
        RECT 54.960 0.180 55.260 0.480 ;
        RECT 55.450 0.180 55.750 0.480 ;
        RECT 55.940 0.180 56.240 0.480 ;
        RECT 58.200 0.180 58.500 0.480 ;
        RECT 58.690 0.180 58.990 0.480 ;
        RECT 59.180 0.180 59.480 0.480 ;
        RECT 59.670 0.180 59.970 0.480 ;
        RECT 60.160 0.180 60.460 0.480 ;
        RECT 60.650 0.180 60.950 0.480 ;
        RECT 61.140 0.180 61.440 0.480 ;
        RECT 61.630 0.180 61.930 0.480 ;
        RECT 63.710 0.180 64.010 0.480 ;
        RECT 64.200 0.180 64.500 0.480 ;
        RECT 64.690 0.180 64.990 0.480 ;
        RECT 65.180 0.180 65.480 0.480 ;
        RECT 65.670 0.180 65.970 0.480 ;
        RECT 66.160 0.180 66.460 0.480 ;
        RECT 66.650 0.180 66.950 0.480 ;
        RECT 67.140 0.180 67.440 0.480 ;
        RECT 69.350 0.180 69.650 0.480 ;
        RECT 69.840 0.180 70.140 0.480 ;
        RECT 70.330 0.180 70.630 0.480 ;
        RECT 70.820 0.180 71.120 0.480 ;
        RECT 72.670 0.180 72.970 0.480 ;
        RECT 73.160 0.180 73.460 0.480 ;
        RECT 73.650 0.180 73.950 0.480 ;
        RECT 75.910 0.180 76.210 0.480 ;
        RECT 76.400 0.180 76.700 0.480 ;
        RECT 76.890 0.180 77.190 0.480 ;
        RECT 77.380 0.180 77.680 0.480 ;
        RECT 77.870 0.180 78.170 0.480 ;
        RECT 78.360 0.180 78.660 0.480 ;
        RECT 78.850 0.180 79.150 0.480 ;
        RECT 79.340 0.180 79.640 0.480 ;
        RECT 81.420 0.180 81.720 0.480 ;
        RECT 81.910 0.180 82.210 0.480 ;
        RECT 82.400 0.180 82.700 0.480 ;
        RECT 82.890 0.180 83.190 0.480 ;
        RECT 83.380 0.180 83.680 0.480 ;
        RECT 83.870 0.180 84.170 0.480 ;
        RECT 84.360 0.180 84.660 0.480 ;
        RECT 84.850 0.180 85.150 0.480 ;
        RECT 87.060 0.180 87.360 0.480 ;
        RECT 87.550 0.180 87.850 0.480 ;
        RECT 88.040 0.180 88.340 0.480 ;
        RECT 88.530 0.180 88.830 0.480 ;
        RECT 90.380 0.180 90.680 0.480 ;
        RECT 90.870 0.180 91.170 0.480 ;
        RECT 91.360 0.180 91.660 0.480 ;
        RECT 93.620 0.180 93.920 0.480 ;
        RECT 94.110 0.180 94.410 0.480 ;
        RECT 94.600 0.180 94.900 0.480 ;
        RECT 95.090 0.180 95.390 0.480 ;
        RECT 95.580 0.180 95.880 0.480 ;
        RECT 96.070 0.180 96.370 0.480 ;
        RECT 96.560 0.180 96.860 0.480 ;
        RECT 97.050 0.180 97.350 0.480 ;
        RECT 99.130 0.180 99.430 0.480 ;
        RECT 99.620 0.180 99.920 0.480 ;
        RECT 100.110 0.180 100.410 0.480 ;
        RECT 100.600 0.180 100.900 0.480 ;
        RECT 101.090 0.180 101.390 0.480 ;
        RECT 101.580 0.180 101.880 0.480 ;
        RECT 102.070 0.180 102.370 0.480 ;
        RECT 102.560 0.180 102.860 0.480 ;
        RECT 104.770 0.180 105.070 0.480 ;
        RECT 105.260 0.180 105.560 0.480 ;
        RECT 105.750 0.180 106.050 0.480 ;
        RECT 106.240 0.180 106.540 0.480 ;
      LAYER met1 ;
        RECT 8.400 29.270 97.550 29.750 ;
        RECT -1.000 25.280 4.565 25.760 ;
        RECT 2.180 24.010 10.340 24.310 ;
        RECT 5.760 23.950 10.340 24.010 ;
        RECT 11.295 23.950 28.050 24.310 ;
        RECT 29.005 23.950 45.760 24.310 ;
        RECT 46.715 23.950 63.470 24.310 ;
        RECT 64.425 23.950 81.180 24.310 ;
        RECT 82.135 23.950 100.220 24.310 ;
        RECT 101.000 24.015 103.005 24.380 ;
        RECT -1.000 22.560 4.565 23.040 ;
        RECT 5.760 17.360 6.120 23.950 ;
        RECT 9.980 22.950 10.340 23.950 ;
        RECT 20.960 22.950 21.320 23.950 ;
        RECT 27.690 22.950 28.050 23.950 ;
        RECT 38.670 22.950 39.030 23.950 ;
        RECT 45.400 22.950 45.760 23.950 ;
        RECT 56.380 22.950 56.740 23.950 ;
        RECT 63.110 22.950 63.470 23.950 ;
        RECT 74.090 22.950 74.450 23.950 ;
        RECT 80.820 22.950 81.180 23.950 ;
        RECT 91.800 22.950 92.160 23.950 ;
        RECT 9.370 22.590 13.640 22.950 ;
        RECT 14.890 22.590 19.160 22.950 ;
        RECT 20.410 22.590 21.910 22.950 ;
        RECT 23.740 22.590 25.240 22.950 ;
        RECT 27.080 22.590 31.350 22.950 ;
        RECT 32.600 22.590 36.870 22.950 ;
        RECT 38.120 22.590 39.620 22.950 ;
        RECT 41.450 22.590 42.950 22.950 ;
        RECT 44.790 22.590 49.060 22.950 ;
        RECT 50.310 22.590 54.580 22.950 ;
        RECT 55.830 22.590 57.330 22.950 ;
        RECT 59.160 22.590 60.660 22.950 ;
        RECT 62.500 22.590 66.770 22.950 ;
        RECT 68.020 22.590 72.290 22.950 ;
        RECT 73.540 22.590 75.040 22.950 ;
        RECT 76.870 22.590 78.370 22.950 ;
        RECT 80.210 22.590 84.480 22.950 ;
        RECT 85.730 22.590 90.000 22.950 ;
        RECT 91.250 22.590 92.750 22.950 ;
        RECT 94.580 22.590 96.080 22.950 ;
        RECT 15.505 21.590 15.865 22.590 ;
        RECT 24.290 21.590 24.650 22.590 ;
        RECT 33.215 21.590 33.575 22.590 ;
        RECT 42.000 21.590 42.360 22.590 ;
        RECT 50.925 21.590 51.285 22.590 ;
        RECT 59.710 21.590 60.070 22.590 ;
        RECT 68.635 21.590 68.995 22.590 ;
        RECT 77.420 21.590 77.780 22.590 ;
        RECT 86.345 21.590 86.705 22.590 ;
        RECT 95.130 21.590 95.490 22.590 ;
        RECT -2.510 17.000 6.120 17.360 ;
        RECT 7.120 21.230 15.865 21.590 ;
        RECT 16.815 21.230 33.575 21.590 ;
        RECT 34.525 21.230 51.285 21.590 ;
        RECT 52.235 21.230 68.995 21.590 ;
        RECT 69.945 21.230 86.705 21.590 ;
        RECT 87.655 21.230 98.860 21.590 ;
        RECT -2.510 5.890 -2.150 17.000 ;
        RECT 7.120 16.000 7.480 21.230 ;
        RECT -1.150 15.640 7.480 16.000 ;
        RECT 8.480 15.670 97.550 16.150 ;
        RECT 98.500 16.000 98.860 21.230 ;
        RECT 99.860 17.360 100.220 23.950 ;
        RECT 102.000 18.500 103.000 19.515 ;
        RECT 107.515 18.500 108.500 19.500 ;
        RECT 99.860 17.000 109.360 17.360 ;
        RECT 98.500 15.640 108.000 16.000 ;
        RECT -1.150 8.610 -0.790 15.640 ;
        RECT 0.000 13.690 106.780 14.170 ;
        RECT 107.640 8.610 108.000 15.640 ;
        RECT -1.150 8.250 9.895 8.610 ;
        RECT 10.845 8.250 27.605 8.610 ;
        RECT 28.555 8.250 45.315 8.610 ;
        RECT 46.265 8.250 63.025 8.610 ;
        RECT 63.975 8.250 80.735 8.610 ;
        RECT 81.685 8.250 98.445 8.610 ;
        RECT 99.395 8.250 108.000 8.610 ;
        RECT 2.060 7.250 2.420 8.250 ;
        RECT 10.845 7.250 11.205 8.250 ;
        RECT 19.770 7.250 20.130 8.250 ;
        RECT 28.555 7.250 28.915 8.250 ;
        RECT 37.480 7.250 37.840 8.250 ;
        RECT 46.265 7.250 46.625 8.250 ;
        RECT 55.190 7.250 55.550 8.250 ;
        RECT 63.975 7.250 64.335 8.250 ;
        RECT 72.900 7.250 73.260 8.250 ;
        RECT 81.685 7.250 82.045 8.250 ;
        RECT 90.610 7.250 90.970 8.250 ;
        RECT 99.395 7.250 99.755 8.250 ;
        RECT 1.470 6.890 2.970 7.250 ;
        RECT 4.800 6.890 6.300 7.250 ;
        RECT 7.550 6.890 11.820 7.250 ;
        RECT 13.070 6.890 17.340 7.250 ;
        RECT 19.180 6.890 20.680 7.250 ;
        RECT 22.510 6.890 24.010 7.250 ;
        RECT 25.260 6.890 29.530 7.250 ;
        RECT 30.780 6.890 35.050 7.250 ;
        RECT 36.890 6.890 38.390 7.250 ;
        RECT 40.220 6.890 41.720 7.250 ;
        RECT 42.970 6.890 47.240 7.250 ;
        RECT 48.490 6.890 52.760 7.250 ;
        RECT 54.600 6.890 56.100 7.250 ;
        RECT 57.930 6.890 59.430 7.250 ;
        RECT 60.680 6.890 64.950 7.250 ;
        RECT 66.200 6.890 70.470 7.250 ;
        RECT 72.310 6.890 73.810 7.250 ;
        RECT 75.640 6.890 77.140 7.250 ;
        RECT 78.390 6.890 82.660 7.250 ;
        RECT 83.910 6.890 88.180 7.250 ;
        RECT 90.020 6.890 91.520 7.250 ;
        RECT 93.350 6.890 94.850 7.250 ;
        RECT 96.100 6.890 100.370 7.250 ;
        RECT 101.620 6.890 105.890 7.250 ;
        RECT 5.390 5.890 5.750 6.890 ;
        RECT 16.370 5.890 16.730 6.890 ;
        RECT 23.100 5.890 23.460 6.890 ;
        RECT 34.080 5.890 34.440 6.890 ;
        RECT 40.810 5.890 41.170 6.890 ;
        RECT 51.790 5.890 52.150 6.890 ;
        RECT 58.520 5.890 58.880 6.890 ;
        RECT 69.500 5.890 69.860 6.890 ;
        RECT 76.230 5.890 76.590 6.890 ;
        RECT 87.210 5.890 87.570 6.890 ;
        RECT 93.940 5.890 94.300 6.890 ;
        RECT 104.920 5.890 105.280 6.890 ;
        RECT 109.000 5.890 109.360 17.000 ;
        RECT -2.510 5.530 15.415 5.890 ;
        RECT 16.370 5.530 33.125 5.890 ;
        RECT 34.080 5.530 50.835 5.890 ;
        RECT 51.790 5.530 68.545 5.890 ;
        RECT 69.500 5.530 86.255 5.890 ;
        RECT 87.210 5.530 103.965 5.890 ;
        RECT 104.920 5.530 109.360 5.890 ;
        RECT 0.000 0.090 106.780 0.570 ;
      LAYER via ;
        RECT 12.000 15.770 12.260 16.030 ;
        RECT 12.370 15.770 12.630 16.030 ;
        RECT 12.740 15.770 13.000 16.030 ;
        RECT 18.000 15.770 18.260 16.030 ;
        RECT 18.370 15.770 18.630 16.030 ;
        RECT 18.740 15.770 19.000 16.030 ;
        RECT 24.000 15.770 24.260 16.030 ;
        RECT 24.370 15.770 24.630 16.030 ;
        RECT 24.740 15.770 25.000 16.030 ;
        RECT 30.000 15.770 30.260 16.030 ;
        RECT 30.370 15.770 30.630 16.030 ;
        RECT 30.740 15.770 31.000 16.030 ;
        RECT 36.000 15.770 36.260 16.030 ;
        RECT 36.370 15.770 36.630 16.030 ;
        RECT 36.740 15.770 37.000 16.030 ;
        RECT 42.000 15.770 42.260 16.030 ;
        RECT 42.370 15.770 42.630 16.030 ;
        RECT 42.740 15.770 43.000 16.030 ;
        RECT 48.000 15.770 48.260 16.030 ;
        RECT 48.370 15.770 48.630 16.030 ;
        RECT 48.740 15.770 49.000 16.030 ;
        RECT 54.000 15.770 54.260 16.030 ;
        RECT 54.370 15.770 54.630 16.030 ;
        RECT 54.740 15.770 55.000 16.030 ;
        RECT 60.000 15.770 60.260 16.030 ;
        RECT 60.370 15.770 60.630 16.030 ;
        RECT 60.740 15.770 61.000 16.030 ;
        RECT 66.000 15.770 66.260 16.030 ;
        RECT 66.370 15.770 66.630 16.030 ;
        RECT 66.740 15.770 67.000 16.030 ;
        RECT 72.000 15.770 72.260 16.030 ;
        RECT 72.370 15.770 72.630 16.030 ;
        RECT 72.740 15.770 73.000 16.030 ;
        RECT 78.000 15.770 78.260 16.030 ;
        RECT 78.370 15.770 78.630 16.030 ;
        RECT 78.740 15.770 79.000 16.030 ;
        RECT 84.000 15.770 84.260 16.030 ;
        RECT 84.370 15.770 84.630 16.030 ;
        RECT 84.740 15.770 85.000 16.030 ;
        RECT 90.000 15.770 90.260 16.030 ;
        RECT 90.370 15.770 90.630 16.030 ;
        RECT 90.740 15.770 91.000 16.030 ;
        RECT 96.000 15.770 96.260 16.030 ;
        RECT 96.370 15.770 96.630 16.030 ;
        RECT 96.740 15.770 97.000 16.030 ;
        RECT 102.070 19.100 102.410 19.440 ;
        RECT 102.590 19.100 102.930 19.440 ;
        RECT 102.070 18.580 102.410 18.920 ;
        RECT 102.590 18.580 102.930 18.920 ;
        RECT 107.585 19.080 107.925 19.420 ;
        RECT 108.075 19.080 108.415 19.420 ;
        RECT 107.585 18.580 107.925 18.920 ;
        RECT 108.075 18.580 108.415 18.920 ;
        RECT 0.000 13.790 0.260 14.050 ;
        RECT 0.370 13.790 0.630 14.050 ;
        RECT 0.740 13.790 1.000 14.050 ;
        RECT 6.000 13.790 6.260 14.050 ;
        RECT 6.370 13.790 6.630 14.050 ;
        RECT 6.740 13.790 7.000 14.050 ;
        RECT 12.000 13.790 12.260 14.050 ;
        RECT 12.370 13.790 12.630 14.050 ;
        RECT 12.740 13.790 13.000 14.050 ;
        RECT 18.000 13.790 18.260 14.050 ;
        RECT 18.370 13.790 18.630 14.050 ;
        RECT 18.740 13.790 19.000 14.050 ;
        RECT 24.000 13.790 24.260 14.050 ;
        RECT 24.370 13.790 24.630 14.050 ;
        RECT 24.740 13.790 25.000 14.050 ;
        RECT 30.000 13.790 30.260 14.050 ;
        RECT 30.370 13.790 30.630 14.050 ;
        RECT 30.740 13.790 31.000 14.050 ;
        RECT 36.000 13.790 36.260 14.050 ;
        RECT 36.370 13.790 36.630 14.050 ;
        RECT 36.740 13.790 37.000 14.050 ;
        RECT 42.000 13.790 42.260 14.050 ;
        RECT 42.370 13.790 42.630 14.050 ;
        RECT 42.740 13.790 43.000 14.050 ;
        RECT 48.000 13.790 48.260 14.050 ;
        RECT 48.370 13.790 48.630 14.050 ;
        RECT 48.740 13.790 49.000 14.050 ;
        RECT 54.000 13.790 54.260 14.050 ;
        RECT 54.370 13.790 54.630 14.050 ;
        RECT 54.740 13.790 55.000 14.050 ;
        RECT 60.000 13.790 60.260 14.050 ;
        RECT 60.370 13.790 60.630 14.050 ;
        RECT 60.740 13.790 61.000 14.050 ;
        RECT 66.000 13.790 66.260 14.050 ;
        RECT 66.370 13.790 66.630 14.050 ;
        RECT 66.740 13.790 67.000 14.050 ;
        RECT 72.000 13.790 72.260 14.050 ;
        RECT 72.370 13.790 72.630 14.050 ;
        RECT 72.740 13.790 73.000 14.050 ;
        RECT 78.000 13.790 78.260 14.050 ;
        RECT 78.370 13.790 78.630 14.050 ;
        RECT 78.740 13.790 79.000 14.050 ;
        RECT 84.000 13.790 84.260 14.050 ;
        RECT 84.370 13.790 84.630 14.050 ;
        RECT 84.740 13.790 85.000 14.050 ;
        RECT 90.000 13.790 90.260 14.050 ;
        RECT 90.370 13.790 90.630 14.050 ;
        RECT 90.740 13.790 91.000 14.050 ;
        RECT 96.000 13.790 96.260 14.050 ;
        RECT 96.370 13.790 96.630 14.050 ;
        RECT 96.740 13.790 97.000 14.050 ;
        RECT 102.000 13.790 102.260 14.050 ;
        RECT 102.370 13.790 102.630 14.050 ;
        RECT 102.740 13.790 103.000 14.050 ;
        RECT 105.780 13.790 106.040 14.050 ;
        RECT 106.150 13.790 106.410 14.050 ;
        RECT 106.520 13.790 106.780 14.050 ;
      LAYER met2 ;
        RECT 102.000 18.500 103.000 19.515 ;
        RECT 107.515 18.500 108.500 19.500 ;
        RECT 12.000 15.700 13.000 16.100 ;
        RECT 18.000 15.700 19.000 16.100 ;
        RECT 24.000 15.700 25.000 16.100 ;
        RECT 30.000 15.700 31.000 16.100 ;
        RECT 36.000 15.700 37.000 16.100 ;
        RECT 42.000 15.700 43.000 16.100 ;
        RECT 48.000 15.700 49.000 16.100 ;
        RECT 54.000 15.700 55.000 16.100 ;
        RECT 60.000 15.700 61.000 16.100 ;
        RECT 66.000 15.700 67.000 16.100 ;
        RECT 72.000 15.700 73.000 16.100 ;
        RECT 78.000 15.700 79.000 16.100 ;
        RECT 84.000 15.700 85.000 16.100 ;
        RECT 90.000 15.700 91.000 16.100 ;
        RECT 96.000 15.700 97.000 16.100 ;
        RECT 0.000 13.720 1.000 14.120 ;
        RECT 6.000 13.720 7.000 14.120 ;
        RECT 12.000 13.720 13.000 14.120 ;
        RECT 18.000 13.720 19.000 14.120 ;
        RECT 24.000 13.720 25.000 14.120 ;
        RECT 30.000 13.720 31.000 14.120 ;
        RECT 36.000 13.720 37.000 14.120 ;
        RECT 42.000 13.720 43.000 14.120 ;
        RECT 48.000 13.720 49.000 14.120 ;
        RECT 54.000 13.720 55.000 14.120 ;
        RECT 60.000 13.720 61.000 14.120 ;
        RECT 66.000 13.720 67.000 14.120 ;
        RECT 72.000 13.720 73.000 14.120 ;
        RECT 78.000 13.720 79.000 14.120 ;
        RECT 84.000 13.720 85.000 14.120 ;
        RECT 90.000 13.720 91.000 14.120 ;
        RECT 96.000 13.720 97.000 14.120 ;
        RECT 102.000 13.720 103.000 14.120 ;
        RECT 105.780 13.720 106.780 14.120 ;
      LAYER via2 ;
        RECT 102.040 19.070 102.440 19.470 ;
        RECT 102.560 19.070 102.960 19.470 ;
        RECT 102.040 18.550 102.440 18.950 ;
        RECT 102.560 18.550 102.960 18.950 ;
        RECT 12.100 15.750 12.400 16.050 ;
        RECT 12.600 15.750 12.900 16.050 ;
        RECT 18.100 15.750 18.400 16.050 ;
        RECT 18.600 15.750 18.900 16.050 ;
        RECT 24.100 15.750 24.400 16.050 ;
        RECT 24.600 15.750 24.900 16.050 ;
        RECT 30.100 15.750 30.400 16.050 ;
        RECT 30.600 15.750 30.900 16.050 ;
        RECT 36.100 15.750 36.400 16.050 ;
        RECT 36.600 15.750 36.900 16.050 ;
        RECT 42.100 15.750 42.400 16.050 ;
        RECT 42.600 15.750 42.900 16.050 ;
        RECT 48.100 15.750 48.400 16.050 ;
        RECT 48.600 15.750 48.900 16.050 ;
        RECT 54.100 15.750 54.400 16.050 ;
        RECT 54.600 15.750 54.900 16.050 ;
        RECT 60.100 15.750 60.400 16.050 ;
        RECT 60.600 15.750 60.900 16.050 ;
        RECT 66.100 15.750 66.400 16.050 ;
        RECT 66.600 15.750 66.900 16.050 ;
        RECT 72.100 15.750 72.400 16.050 ;
        RECT 72.600 15.750 72.900 16.050 ;
        RECT 78.100 15.750 78.400 16.050 ;
        RECT 78.600 15.750 78.900 16.050 ;
        RECT 84.100 15.750 84.400 16.050 ;
        RECT 84.600 15.750 84.900 16.050 ;
        RECT 90.100 15.750 90.400 16.050 ;
        RECT 90.600 15.750 90.900 16.050 ;
        RECT 96.100 15.750 96.400 16.050 ;
        RECT 96.600 15.750 96.900 16.050 ;
        RECT 0.100 13.770 0.400 14.070 ;
        RECT 0.600 13.770 0.900 14.070 ;
        RECT 6.100 13.770 6.400 14.070 ;
        RECT 6.600 13.770 6.900 14.070 ;
        RECT 12.100 13.770 12.400 14.070 ;
        RECT 12.600 13.770 12.900 14.070 ;
        RECT 18.100 13.770 18.400 14.070 ;
        RECT 18.600 13.770 18.900 14.070 ;
        RECT 24.100 13.770 24.400 14.070 ;
        RECT 24.600 13.770 24.900 14.070 ;
        RECT 30.100 13.770 30.400 14.070 ;
        RECT 30.600 13.770 30.900 14.070 ;
        RECT 36.100 13.770 36.400 14.070 ;
        RECT 36.600 13.770 36.900 14.070 ;
        RECT 42.100 13.770 42.400 14.070 ;
        RECT 42.600 13.770 42.900 14.070 ;
        RECT 48.100 13.770 48.400 14.070 ;
        RECT 48.600 13.770 48.900 14.070 ;
        RECT 54.100 13.770 54.400 14.070 ;
        RECT 54.600 13.770 54.900 14.070 ;
        RECT 60.100 13.770 60.400 14.070 ;
        RECT 60.600 13.770 60.900 14.070 ;
        RECT 66.100 13.770 66.400 14.070 ;
        RECT 66.600 13.770 66.900 14.070 ;
        RECT 72.100 13.770 72.400 14.070 ;
        RECT 72.600 13.770 72.900 14.070 ;
        RECT 78.100 13.770 78.400 14.070 ;
        RECT 78.600 13.770 78.900 14.070 ;
        RECT 84.100 13.770 84.400 14.070 ;
        RECT 84.600 13.770 84.900 14.070 ;
        RECT 90.100 13.770 90.400 14.070 ;
        RECT 90.600 13.770 90.900 14.070 ;
        RECT 96.100 13.770 96.400 14.070 ;
        RECT 96.600 13.770 96.900 14.070 ;
        RECT 102.100 13.770 102.400 14.070 ;
        RECT 102.600 13.770 102.900 14.070 ;
        RECT 105.880 13.770 106.180 14.070 ;
        RECT 106.380 13.770 106.680 14.070 ;
      LAYER met3 ;
        RECT 12.000 15.670 13.000 16.150 ;
        RECT 18.000 15.670 19.000 16.150 ;
        RECT 24.000 15.670 25.000 16.150 ;
        RECT 30.000 15.670 31.000 16.150 ;
        RECT 36.000 15.670 37.000 16.150 ;
        RECT 42.000 15.670 43.000 16.150 ;
        RECT 48.000 15.670 49.000 16.150 ;
        RECT 54.000 15.670 55.000 16.150 ;
        RECT 60.000 15.670 61.000 16.150 ;
        RECT 66.000 15.670 67.000 16.150 ;
        RECT 72.000 15.670 73.000 16.150 ;
        RECT 78.000 15.670 79.000 16.150 ;
        RECT 84.000 15.670 85.000 16.150 ;
        RECT 90.000 15.670 91.000 16.150 ;
        RECT 96.000 15.670 97.000 16.150 ;
        RECT 102.000 15.670 103.000 19.515 ;
        RECT 0.000 14.170 106.780 15.670 ;
        RECT 0.000 13.690 1.000 14.170 ;
        RECT 6.000 13.690 7.000 14.170 ;
        RECT 12.000 13.690 13.000 14.170 ;
        RECT 18.000 13.690 19.000 14.170 ;
        RECT 24.000 13.690 25.000 14.170 ;
        RECT 30.000 13.690 31.000 14.170 ;
        RECT 36.000 13.690 37.000 14.170 ;
        RECT 42.000 13.690 43.000 14.170 ;
        RECT 48.000 13.690 49.000 14.170 ;
        RECT 54.000 13.690 55.000 14.170 ;
        RECT 60.000 13.690 61.000 14.170 ;
        RECT 66.000 13.690 67.000 14.170 ;
        RECT 72.000 13.690 73.000 14.170 ;
        RECT 78.000 13.690 79.000 14.170 ;
        RECT 84.000 13.690 85.000 14.170 ;
        RECT 90.000 13.690 91.000 14.170 ;
        RECT 96.000 13.690 97.000 14.170 ;
        RECT 102.000 13.690 103.000 14.170 ;
        RECT 105.780 13.690 106.780 14.170 ;
  END
END ring_osc
MACRO vco_w6_r100
  CLASS BLOCK ;
  FOREIGN vco_w6_r100 ;
  ORIGIN 5.000 38.000 ;
  SIZE 122.000 BY 105.000 ;
  SYMMETRY X Y R90 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 87.420 7.250 87.800 7.300 ;
        RECT 86.470 6.890 87.800 7.250 ;
        RECT 87.420 6.840 87.800 6.890 ;
        RECT 89.290 7.250 89.670 7.300 ;
        RECT 89.290 6.890 90.620 7.250 ;
        RECT 89.290 6.840 89.670 6.890 ;
        RECT 91.730 0.750 92.030 13.340 ;
        RECT 95.960 7.250 96.340 7.300 ;
        RECT 95.960 6.890 97.290 7.250 ;
        RECT 95.960 6.840 96.340 6.890 ;
        RECT 106.105 0.750 106.405 13.340 ;
      LAYER mcon ;
        RECT 86.470 6.920 86.770 7.220 ;
        RECT 86.960 6.920 87.260 7.220 ;
        RECT 87.450 6.920 87.750 7.220 ;
        RECT 89.340 6.920 89.640 7.220 ;
        RECT 89.830 6.920 90.130 7.220 ;
        RECT 90.320 6.920 90.620 7.220 ;
        RECT 96.010 6.920 96.310 7.220 ;
        RECT 96.500 6.920 96.800 7.220 ;
        RECT 96.990 6.920 97.290 7.220 ;
        RECT 91.730 5.560 92.030 5.860 ;
        RECT 106.105 5.560 106.405 5.860 ;
      LAYER met1 ;
        RECT 86.410 6.890 90.680 7.250 ;
        RECT 95.850 6.890 97.350 7.250 ;
        RECT 89.710 5.890 90.070 6.890 ;
        RECT 96.440 5.890 96.800 6.890 ;
        RECT 89.710 5.530 106.465 5.890 ;
      LAYER via ;
        RECT 91.140 5.530 91.500 5.890 ;
      LAYER met2 ;
        RECT 91.110 -38.420 91.530 5.890 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 69.710 7.250 70.090 7.300 ;
        RECT 68.760 6.890 70.090 7.250 ;
        RECT 69.710 6.840 70.090 6.890 ;
        RECT 71.580 7.250 71.960 7.300 ;
        RECT 71.580 6.890 72.910 7.250 ;
        RECT 71.580 6.840 71.960 6.890 ;
        RECT 74.020 0.750 74.320 13.340 ;
        RECT 78.250 7.250 78.630 7.300 ;
        RECT 78.250 6.890 79.580 7.250 ;
        RECT 78.250 6.840 78.630 6.890 ;
        RECT 88.395 0.750 88.695 13.340 ;
      LAYER mcon ;
        RECT 68.760 6.920 69.060 7.220 ;
        RECT 69.250 6.920 69.550 7.220 ;
        RECT 69.740 6.920 70.040 7.220 ;
        RECT 71.630 6.920 71.930 7.220 ;
        RECT 72.120 6.920 72.420 7.220 ;
        RECT 72.610 6.920 72.910 7.220 ;
        RECT 78.300 6.920 78.600 7.220 ;
        RECT 78.790 6.920 79.090 7.220 ;
        RECT 79.280 6.920 79.580 7.220 ;
        RECT 74.020 5.560 74.320 5.860 ;
        RECT 88.395 5.560 88.695 5.860 ;
      LAYER met1 ;
        RECT 68.700 6.890 72.970 7.250 ;
        RECT 78.140 6.890 79.640 7.250 ;
        RECT 72.000 5.890 72.360 6.890 ;
        RECT 78.730 5.890 79.090 6.890 ;
        RECT 72.000 5.530 88.755 5.890 ;
      LAYER via ;
        RECT 74.340 5.530 74.700 5.890 ;
      LAYER met2 ;
        RECT 74.310 -38.420 74.730 5.890 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 52.000 7.250 52.380 7.300 ;
        RECT 51.050 6.890 52.380 7.250 ;
        RECT 52.000 6.840 52.380 6.890 ;
        RECT 53.870 7.250 54.250 7.300 ;
        RECT 53.870 6.890 55.200 7.250 ;
        RECT 53.870 6.840 54.250 6.890 ;
        RECT 56.310 0.750 56.610 13.340 ;
        RECT 60.540 7.250 60.920 7.300 ;
        RECT 60.540 6.890 61.870 7.250 ;
        RECT 60.540 6.840 60.920 6.890 ;
        RECT 70.685 0.750 70.985 13.340 ;
      LAYER mcon ;
        RECT 51.050 6.920 51.350 7.220 ;
        RECT 51.540 6.920 51.840 7.220 ;
        RECT 52.030 6.920 52.330 7.220 ;
        RECT 53.920 6.920 54.220 7.220 ;
        RECT 54.410 6.920 54.710 7.220 ;
        RECT 54.900 6.920 55.200 7.220 ;
        RECT 60.590 6.920 60.890 7.220 ;
        RECT 61.080 6.920 61.380 7.220 ;
        RECT 61.570 6.920 61.870 7.220 ;
        RECT 56.310 5.560 56.610 5.860 ;
        RECT 70.685 5.560 70.985 5.860 ;
      LAYER met1 ;
        RECT 50.990 6.890 55.260 7.250 ;
        RECT 60.430 6.890 61.930 7.250 ;
        RECT 54.290 5.890 54.650 6.890 ;
        RECT 61.020 5.890 61.380 6.890 ;
        RECT 54.290 5.530 71.045 5.890 ;
      LAYER via ;
        RECT 61.020 5.530 61.380 5.890 ;
      LAYER met2 ;
        RECT 60.990 -38.420 61.410 5.890 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 34.290 7.250 34.670 7.300 ;
        RECT 33.340 6.890 34.670 7.250 ;
        RECT 34.290 6.840 34.670 6.890 ;
        RECT 36.160 7.250 36.540 7.300 ;
        RECT 36.160 6.890 37.490 7.250 ;
        RECT 36.160 6.840 36.540 6.890 ;
        RECT 38.600 0.750 38.900 13.340 ;
        RECT 42.830 7.250 43.210 7.300 ;
        RECT 42.830 6.890 44.160 7.250 ;
        RECT 42.830 6.840 43.210 6.890 ;
        RECT 52.975 0.750 53.275 13.340 ;
      LAYER mcon ;
        RECT 33.340 6.920 33.640 7.220 ;
        RECT 33.830 6.920 34.130 7.220 ;
        RECT 34.320 6.920 34.620 7.220 ;
        RECT 36.210 6.920 36.510 7.220 ;
        RECT 36.700 6.920 37.000 7.220 ;
        RECT 37.190 6.920 37.490 7.220 ;
        RECT 42.880 6.920 43.180 7.220 ;
        RECT 43.370 6.920 43.670 7.220 ;
        RECT 43.860 6.920 44.160 7.220 ;
        RECT 38.600 5.560 38.900 5.860 ;
        RECT 52.975 5.560 53.275 5.860 ;
      LAYER met1 ;
        RECT 33.280 6.890 37.550 7.250 ;
        RECT 42.720 6.890 44.220 7.250 ;
        RECT 36.580 5.890 36.940 6.890 ;
        RECT 43.310 5.890 43.670 6.890 ;
        RECT 36.580 5.530 53.335 5.890 ;
      LAYER via ;
        RECT 38.030 5.530 38.390 5.890 ;
      LAYER met2 ;
        RECT 38.000 -38.420 38.420 5.890 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 16.580 7.250 16.960 7.300 ;
        RECT 15.630 6.890 16.960 7.250 ;
        RECT 16.580 6.840 16.960 6.890 ;
        RECT 18.450 7.250 18.830 7.300 ;
        RECT 18.450 6.890 19.780 7.250 ;
        RECT 18.450 6.840 18.830 6.890 ;
        RECT 20.890 0.750 21.190 13.340 ;
        RECT 25.120 7.250 25.500 7.300 ;
        RECT 25.120 6.890 26.450 7.250 ;
        RECT 25.120 6.840 25.500 6.890 ;
        RECT 35.265 0.750 35.565 13.340 ;
      LAYER mcon ;
        RECT 15.630 6.920 15.930 7.220 ;
        RECT 16.120 6.920 16.420 7.220 ;
        RECT 16.610 6.920 16.910 7.220 ;
        RECT 18.500 6.920 18.800 7.220 ;
        RECT 18.990 6.920 19.290 7.220 ;
        RECT 19.480 6.920 19.780 7.220 ;
        RECT 25.170 6.920 25.470 7.220 ;
        RECT 25.660 6.920 25.960 7.220 ;
        RECT 26.150 6.920 26.450 7.220 ;
        RECT 20.890 5.560 21.190 5.860 ;
        RECT 35.265 5.560 35.565 5.860 ;
      LAYER met1 ;
        RECT 15.570 6.890 19.840 7.250 ;
        RECT 25.010 6.890 26.510 7.250 ;
        RECT 18.870 5.890 19.230 6.890 ;
        RECT 25.600 5.890 25.960 6.890 ;
        RECT 18.870 5.530 35.625 5.890 ;
      LAYER via ;
        RECT 20.280 5.530 20.640 5.890 ;
      LAYER met2 ;
        RECT 20.250 -38.420 20.670 5.890 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 6.245500 ;
    PORT
      LAYER li1 ;
        RECT 3.310 24.925 3.905 25.265 ;
        RECT 3.310 23.605 3.485 24.925 ;
        RECT 3.310 23.480 3.905 23.605 ;
        RECT 4.710 23.480 5.010 24.310 ;
        RECT 3.310 23.180 5.010 23.480 ;
        RECT 3.310 23.055 3.905 23.180 ;
        RECT 12.880 22.950 13.260 23.000 ;
        RECT 11.930 22.590 13.260 22.950 ;
        RECT 12.880 22.540 13.260 22.590 ;
        RECT 14.750 22.950 15.130 23.000 ;
        RECT 14.750 22.590 16.080 22.950 ;
        RECT 14.750 22.540 15.130 22.590 ;
        RECT 3.180 0.750 3.480 13.340 ;
        RECT 7.410 7.250 7.790 7.300 ;
        RECT 7.410 6.890 8.740 7.250 ;
        RECT 7.410 6.840 7.790 6.890 ;
        RECT 17.555 0.750 17.855 13.340 ;
      LAYER mcon ;
        RECT 4.740 24.040 4.980 24.280 ;
        RECT 11.930 22.620 12.230 22.920 ;
        RECT 12.420 22.620 12.720 22.920 ;
        RECT 12.910 22.620 13.210 22.920 ;
        RECT 14.800 22.620 15.100 22.920 ;
        RECT 15.290 22.620 15.590 22.920 ;
        RECT 15.780 22.620 16.080 22.920 ;
        RECT 7.460 6.920 7.760 7.220 ;
        RECT 7.950 6.920 8.250 7.220 ;
        RECT 8.440 6.920 8.740 7.220 ;
        RECT 3.180 5.560 3.480 5.860 ;
        RECT 17.555 5.560 17.855 5.860 ;
      LAYER met1 ;
        RECT 4.680 24.010 12.840 24.310 ;
        RECT 8.260 23.950 12.840 24.010 ;
        RECT 8.260 17.360 8.620 23.950 ;
        RECT 12.480 22.950 12.840 23.950 ;
        RECT 11.870 22.590 16.140 22.950 ;
        RECT -0.010 17.000 8.620 17.360 ;
        RECT -0.010 5.890 0.350 17.000 ;
        RECT 7.300 6.890 8.800 7.250 ;
        RECT 7.890 5.890 8.250 6.890 ;
        RECT -0.010 5.530 17.915 5.890 ;
      LAYER via ;
        RECT 2.140 5.530 2.500 5.890 ;
      LAYER met2 ;
        RECT 2.110 -38.420 2.530 5.890 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 13.855 16.500 14.155 29.090 ;
        RECT 23.920 22.950 24.300 23.000 ;
        RECT 22.970 22.590 24.300 22.950 ;
        RECT 23.920 22.540 24.300 22.590 ;
        RECT 28.230 16.500 28.530 29.090 ;
        RECT 30.590 22.950 30.970 23.000 ;
        RECT 29.640 22.590 30.970 22.950 ;
        RECT 30.590 22.540 30.970 22.590 ;
        RECT 32.460 22.950 32.840 23.000 ;
        RECT 32.460 22.590 33.790 22.950 ;
        RECT 32.460 22.540 32.840 22.590 ;
      LAYER mcon ;
        RECT 13.855 23.980 14.155 24.280 ;
        RECT 28.230 23.980 28.530 24.280 ;
        RECT 22.970 22.620 23.270 22.920 ;
        RECT 23.460 22.620 23.760 22.920 ;
        RECT 23.950 22.620 24.250 22.920 ;
        RECT 29.640 22.620 29.940 22.920 ;
        RECT 30.130 22.620 30.430 22.920 ;
        RECT 30.620 22.620 30.920 22.920 ;
        RECT 32.510 22.620 32.810 22.920 ;
        RECT 33.000 22.620 33.300 22.920 ;
        RECT 33.490 22.620 33.790 22.920 ;
      LAYER met1 ;
        RECT 13.795 23.950 30.550 24.310 ;
        RECT 23.460 22.950 23.820 23.950 ;
        RECT 30.190 22.950 30.550 23.950 ;
        RECT 22.910 22.590 24.410 22.950 ;
        RECT 29.580 22.590 33.850 22.950 ;
      LAYER via ;
        RECT 22.110 23.950 22.470 24.310 ;
      LAYER met2 ;
        RECT 22.080 23.950 22.500 67.420 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 31.565 16.500 31.865 29.090 ;
        RECT 41.630 22.950 42.010 23.000 ;
        RECT 40.680 22.590 42.010 22.950 ;
        RECT 41.630 22.540 42.010 22.590 ;
        RECT 45.940 16.500 46.240 29.090 ;
        RECT 48.300 22.950 48.680 23.000 ;
        RECT 47.350 22.590 48.680 22.950 ;
        RECT 48.300 22.540 48.680 22.590 ;
        RECT 50.170 22.950 50.550 23.000 ;
        RECT 50.170 22.590 51.500 22.950 ;
        RECT 50.170 22.540 50.550 22.590 ;
      LAYER mcon ;
        RECT 31.565 23.980 31.865 24.280 ;
        RECT 45.940 23.980 46.240 24.280 ;
        RECT 40.680 22.620 40.980 22.920 ;
        RECT 41.170 22.620 41.470 22.920 ;
        RECT 41.660 22.620 41.960 22.920 ;
        RECT 47.350 22.620 47.650 22.920 ;
        RECT 47.840 22.620 48.140 22.920 ;
        RECT 48.330 22.620 48.630 22.920 ;
        RECT 50.220 22.620 50.520 22.920 ;
        RECT 50.710 22.620 51.010 22.920 ;
        RECT 51.200 22.620 51.500 22.920 ;
      LAYER met1 ;
        RECT 31.505 23.950 48.260 24.310 ;
        RECT 41.170 22.950 41.530 23.950 ;
        RECT 47.900 22.950 48.260 23.950 ;
        RECT 40.620 22.590 42.120 22.950 ;
        RECT 47.290 22.590 51.560 22.950 ;
      LAYER via ;
        RECT 46.480 23.950 46.840 24.310 ;
      LAYER met2 ;
        RECT 46.450 23.950 46.870 67.420 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 49.275 16.500 49.575 29.090 ;
        RECT 59.340 22.950 59.720 23.000 ;
        RECT 58.390 22.590 59.720 22.950 ;
        RECT 59.340 22.540 59.720 22.590 ;
        RECT 63.650 16.500 63.950 29.090 ;
        RECT 66.010 22.950 66.390 23.000 ;
        RECT 65.060 22.590 66.390 22.950 ;
        RECT 66.010 22.540 66.390 22.590 ;
        RECT 67.880 22.950 68.260 23.000 ;
        RECT 67.880 22.590 69.210 22.950 ;
        RECT 67.880 22.540 68.260 22.590 ;
      LAYER mcon ;
        RECT 49.275 23.980 49.575 24.280 ;
        RECT 63.650 23.980 63.950 24.280 ;
        RECT 58.390 22.620 58.690 22.920 ;
        RECT 58.880 22.620 59.180 22.920 ;
        RECT 59.370 22.620 59.670 22.920 ;
        RECT 65.060 22.620 65.360 22.920 ;
        RECT 65.550 22.620 65.850 22.920 ;
        RECT 66.040 22.620 66.340 22.920 ;
        RECT 67.930 22.620 68.230 22.920 ;
        RECT 68.420 22.620 68.720 22.920 ;
        RECT 68.910 22.620 69.210 22.920 ;
      LAYER met1 ;
        RECT 49.215 23.950 65.970 24.310 ;
        RECT 58.880 22.950 59.240 23.950 ;
        RECT 65.610 22.950 65.970 23.950 ;
        RECT 58.330 22.590 59.830 22.950 ;
        RECT 65.000 22.590 69.270 22.950 ;
      LAYER via ;
        RECT 63.270 23.950 63.630 24.310 ;
      LAYER met2 ;
        RECT 63.240 23.950 63.660 67.420 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 66.985 16.500 67.285 29.090 ;
        RECT 77.050 22.950 77.430 23.000 ;
        RECT 76.100 22.590 77.430 22.950 ;
        RECT 77.050 22.540 77.430 22.590 ;
        RECT 81.360 16.500 81.660 29.090 ;
        RECT 83.720 22.950 84.100 23.000 ;
        RECT 82.770 22.590 84.100 22.950 ;
        RECT 83.720 22.540 84.100 22.590 ;
        RECT 85.590 22.950 85.970 23.000 ;
        RECT 85.590 22.590 86.920 22.950 ;
        RECT 85.590 22.540 85.970 22.590 ;
      LAYER mcon ;
        RECT 66.985 23.980 67.285 24.280 ;
        RECT 81.360 23.980 81.660 24.280 ;
        RECT 76.100 22.620 76.400 22.920 ;
        RECT 76.590 22.620 76.890 22.920 ;
        RECT 77.080 22.620 77.380 22.920 ;
        RECT 82.770 22.620 83.070 22.920 ;
        RECT 83.260 22.620 83.560 22.920 ;
        RECT 83.750 22.620 84.050 22.920 ;
        RECT 85.640 22.620 85.940 22.920 ;
        RECT 86.130 22.620 86.430 22.920 ;
        RECT 86.620 22.620 86.920 22.920 ;
      LAYER met1 ;
        RECT 66.925 23.950 83.680 24.310 ;
        RECT 76.590 22.950 76.950 23.950 ;
        RECT 83.320 22.950 83.680 23.950 ;
        RECT 76.040 22.590 77.540 22.950 ;
        RECT 82.710 22.590 86.980 22.950 ;
      LAYER via ;
        RECT 78.570 23.950 78.930 24.310 ;
      LAYER met2 ;
        RECT 78.540 23.950 78.960 67.420 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 84.695 16.500 84.995 29.090 ;
        RECT 94.760 22.950 95.140 23.000 ;
        RECT 93.810 22.590 95.140 22.950 ;
        RECT 94.760 22.540 95.140 22.590 ;
        RECT 99.070 16.500 99.370 29.090 ;
        RECT 105.130 7.250 105.510 7.300 ;
        RECT 104.180 6.890 105.510 7.250 ;
        RECT 105.130 6.840 105.510 6.890 ;
        RECT 107.000 7.250 107.380 7.300 ;
        RECT 107.000 6.890 108.330 7.250 ;
        RECT 107.000 6.840 107.380 6.890 ;
      LAYER mcon ;
        RECT 84.695 23.980 84.995 24.280 ;
        RECT 99.070 23.980 99.370 24.280 ;
        RECT 93.810 22.620 94.110 22.920 ;
        RECT 94.300 22.620 94.600 22.920 ;
        RECT 94.790 22.620 95.090 22.920 ;
        RECT 104.180 6.920 104.480 7.220 ;
        RECT 104.670 6.920 104.970 7.220 ;
        RECT 105.160 6.920 105.460 7.220 ;
        RECT 107.050 6.920 107.350 7.220 ;
        RECT 107.540 6.920 107.840 7.220 ;
        RECT 108.030 6.920 108.330 7.220 ;
      LAYER met1 ;
        RECT 84.635 23.950 102.720 24.310 ;
        RECT 94.300 22.950 94.660 23.950 ;
        RECT 93.750 22.590 95.250 22.950 ;
        RECT 102.360 17.360 102.720 23.950 ;
        RECT 102.360 17.000 111.860 17.360 ;
        RECT 104.120 6.890 108.390 7.250 ;
        RECT 107.420 5.890 107.780 6.890 ;
        RECT 111.500 5.890 111.860 17.000 ;
        RECT 107.420 5.530 111.860 5.890 ;
      LAYER via ;
        RECT 101.000 23.950 101.360 24.310 ;
      LAYER met2 ;
        RECT 100.970 23.950 101.390 67.420 ;
    END
  END p[10]
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 1.775 24.300 2.235 24.525 ;
        RECT -5.400 24.000 2.235 24.300 ;
        RECT 1.775 23.795 2.235 24.000 ;
      LAYER mcon ;
        RECT -5.380 24.020 -5.120 24.280 ;
      LAYER met1 ;
        RECT -5.450 23.950 -5.050 24.350 ;
    END
  END enb
  PIN input_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 110.015 18.500 111.000 19.500 ;
        RECT 110.015 17.500 110.380 18.500 ;
      LAYER mcon ;
        RECT 110.105 19.100 110.405 19.400 ;
        RECT 110.595 19.100 110.895 19.400 ;
        RECT 110.105 18.600 110.405 18.900 ;
        RECT 110.595 18.600 110.895 18.900 ;
      LAYER met1 ;
        RECT 110.015 18.500 111.000 19.500 ;
      LAYER via ;
        RECT 110.085 19.080 110.425 19.420 ;
        RECT 110.575 19.080 110.915 19.420 ;
        RECT 110.085 18.580 110.425 18.920 ;
        RECT 110.575 18.580 110.915 18.920 ;
      LAYER met2 ;
        RECT 110.010 19.000 118.100 19.500 ;
        RECT 110.015 18.500 111.000 19.000 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.500 24.105 4.180 25.950 ;
        RECT 10.980 22.965 100.050 29.840 ;
        RECT 22.020 22.960 29.210 22.965 ;
        RECT 39.730 22.960 46.920 22.965 ;
        RECT 57.440 22.960 64.630 22.965 ;
        RECT 75.150 22.960 82.340 22.965 ;
        RECT 92.860 22.960 100.050 22.965 ;
        RECT 2.500 6.875 9.690 6.880 ;
        RECT 20.210 6.875 27.400 6.880 ;
        RECT 37.920 6.875 45.110 6.880 ;
        RECT 55.630 6.875 62.820 6.880 ;
        RECT 73.340 6.875 80.530 6.880 ;
        RECT 91.050 6.875 98.240 6.880 ;
        RECT 2.500 0.000 109.280 6.875 ;
      LAYER li1 ;
        RECT 11.160 29.660 13.050 29.690 ;
        RECT 14.840 29.660 18.690 29.690 ;
        RECT 20.350 29.660 24.200 29.690 ;
        RECT 26.040 29.660 27.440 29.690 ;
        RECT 28.870 29.660 30.760 29.690 ;
        RECT 32.550 29.660 36.400 29.690 ;
        RECT 38.060 29.660 41.910 29.690 ;
        RECT 43.750 29.660 45.150 29.690 ;
        RECT 46.580 29.660 48.470 29.690 ;
        RECT 50.260 29.660 54.110 29.690 ;
        RECT 55.770 29.660 59.620 29.690 ;
        RECT 61.460 29.660 62.860 29.690 ;
        RECT 64.290 29.660 66.180 29.690 ;
        RECT 67.970 29.660 71.820 29.690 ;
        RECT 73.480 29.660 77.330 29.690 ;
        RECT 79.170 29.660 80.570 29.690 ;
        RECT 82.000 29.660 83.890 29.690 ;
        RECT 85.680 29.660 89.530 29.690 ;
        RECT 91.190 29.660 95.040 29.690 ;
        RECT 96.880 29.660 98.280 29.690 ;
        RECT 11.160 29.490 99.870 29.660 ;
        RECT 11.160 29.330 13.050 29.490 ;
        RECT 14.840 29.330 18.690 29.490 ;
        RECT 20.350 29.330 24.200 29.490 ;
        RECT 26.040 29.330 27.440 29.490 ;
        RECT 28.870 29.330 30.760 29.490 ;
        RECT 32.550 29.330 36.400 29.490 ;
        RECT 38.060 29.330 41.910 29.490 ;
        RECT 43.750 29.330 45.150 29.490 ;
        RECT 46.580 29.330 48.470 29.490 ;
        RECT 50.260 29.330 54.110 29.490 ;
        RECT 55.770 29.330 59.620 29.490 ;
        RECT 61.460 29.330 62.860 29.490 ;
        RECT 64.290 29.330 66.180 29.490 ;
        RECT 67.970 29.330 71.820 29.490 ;
        RECT 73.480 29.330 77.330 29.490 ;
        RECT 79.170 29.330 80.570 29.490 ;
        RECT 82.000 29.330 83.890 29.490 ;
        RECT 85.680 29.330 89.530 29.490 ;
        RECT 91.190 29.330 95.040 29.490 ;
        RECT 96.880 29.330 98.280 29.490 ;
        RECT 1.690 25.605 2.690 25.770 ;
        RECT 1.690 25.435 3.990 25.605 ;
        RECT 5.685 25.435 7.065 25.605 ;
        RECT 2.205 25.035 3.140 25.435 ;
        RECT 5.960 24.710 6.290 25.435 ;
        RECT 11.160 24.460 11.330 29.330 ;
        RECT 11.670 24.040 11.960 29.330 ;
        RECT 16.050 24.040 16.340 29.330 ;
        RECT 16.680 24.460 16.850 29.330 ;
        RECT 17.190 24.040 17.480 29.330 ;
        RECT 21.570 24.040 21.860 29.330 ;
        RECT 22.200 24.460 22.370 29.330 ;
        RECT 22.710 24.030 23.000 29.330 ;
        RECT 26.040 24.030 26.330 29.330 ;
        RECT 28.870 24.460 29.040 29.330 ;
        RECT 29.380 24.040 29.670 29.330 ;
        RECT 33.760 24.040 34.050 29.330 ;
        RECT 34.390 24.460 34.560 29.330 ;
        RECT 34.900 24.040 35.190 29.330 ;
        RECT 39.280 24.040 39.570 29.330 ;
        RECT 39.910 24.460 40.080 29.330 ;
        RECT 40.420 24.030 40.710 29.330 ;
        RECT 43.750 24.030 44.040 29.330 ;
        RECT 46.580 24.460 46.750 29.330 ;
        RECT 47.090 24.040 47.380 29.330 ;
        RECT 51.470 24.040 51.760 29.330 ;
        RECT 52.100 24.460 52.270 29.330 ;
        RECT 52.610 24.040 52.900 29.330 ;
        RECT 56.990 24.040 57.280 29.330 ;
        RECT 57.620 24.460 57.790 29.330 ;
        RECT 58.130 24.030 58.420 29.330 ;
        RECT 61.460 24.030 61.750 29.330 ;
        RECT 64.290 24.460 64.460 29.330 ;
        RECT 64.800 24.040 65.090 29.330 ;
        RECT 69.180 24.040 69.470 29.330 ;
        RECT 69.810 24.460 69.980 29.330 ;
        RECT 70.320 24.040 70.610 29.330 ;
        RECT 74.700 24.040 74.990 29.330 ;
        RECT 75.330 24.460 75.500 29.330 ;
        RECT 75.840 24.030 76.130 29.330 ;
        RECT 79.170 24.030 79.460 29.330 ;
        RECT 82.000 24.460 82.170 29.330 ;
        RECT 82.510 24.040 82.800 29.330 ;
        RECT 86.890 24.040 87.180 29.330 ;
        RECT 87.520 24.460 87.690 29.330 ;
        RECT 88.030 24.040 88.320 29.330 ;
        RECT 92.410 24.040 92.700 29.330 ;
        RECT 93.040 24.460 93.210 29.330 ;
        RECT 93.550 24.030 93.840 29.330 ;
        RECT 96.880 24.030 97.170 29.330 ;
        RECT 5.380 0.510 5.670 5.810 ;
        RECT 8.710 0.510 9.000 5.810 ;
        RECT 9.340 0.510 9.510 5.380 ;
        RECT 9.850 0.510 10.140 5.800 ;
        RECT 14.230 0.510 14.520 5.800 ;
        RECT 14.860 0.510 15.030 5.380 ;
        RECT 15.370 0.510 15.660 5.800 ;
        RECT 19.750 0.510 20.040 5.800 ;
        RECT 20.380 0.510 20.550 5.380 ;
        RECT 23.090 0.510 23.380 5.810 ;
        RECT 26.420 0.510 26.710 5.810 ;
        RECT 27.050 0.510 27.220 5.380 ;
        RECT 27.560 0.510 27.850 5.800 ;
        RECT 31.940 0.510 32.230 5.800 ;
        RECT 32.570 0.510 32.740 5.380 ;
        RECT 33.080 0.510 33.370 5.800 ;
        RECT 37.460 0.510 37.750 5.800 ;
        RECT 38.090 0.510 38.260 5.380 ;
        RECT 40.800 0.510 41.090 5.810 ;
        RECT 44.130 0.510 44.420 5.810 ;
        RECT 44.760 0.510 44.930 5.380 ;
        RECT 45.270 0.510 45.560 5.800 ;
        RECT 49.650 0.510 49.940 5.800 ;
        RECT 50.280 0.510 50.450 5.380 ;
        RECT 50.790 0.510 51.080 5.800 ;
        RECT 55.170 0.510 55.460 5.800 ;
        RECT 55.800 0.510 55.970 5.380 ;
        RECT 58.510 0.510 58.800 5.810 ;
        RECT 61.840 0.510 62.130 5.810 ;
        RECT 62.470 0.510 62.640 5.380 ;
        RECT 62.980 0.510 63.270 5.800 ;
        RECT 67.360 0.510 67.650 5.800 ;
        RECT 67.990 0.510 68.160 5.380 ;
        RECT 68.500 0.510 68.790 5.800 ;
        RECT 72.880 0.510 73.170 5.800 ;
        RECT 73.510 0.510 73.680 5.380 ;
        RECT 76.220 0.510 76.510 5.810 ;
        RECT 79.550 0.510 79.840 5.810 ;
        RECT 80.180 0.510 80.350 5.380 ;
        RECT 80.690 0.510 80.980 5.800 ;
        RECT 85.070 0.510 85.360 5.800 ;
        RECT 85.700 0.510 85.870 5.380 ;
        RECT 86.210 0.510 86.500 5.800 ;
        RECT 90.590 0.510 90.880 5.800 ;
        RECT 91.220 0.510 91.390 5.380 ;
        RECT 93.930 0.510 94.220 5.810 ;
        RECT 97.260 0.510 97.550 5.810 ;
        RECT 97.890 0.510 98.060 5.380 ;
        RECT 98.400 0.510 98.690 5.800 ;
        RECT 102.780 0.510 103.070 5.800 ;
        RECT 103.410 0.510 103.580 5.380 ;
        RECT 103.920 0.510 104.210 5.800 ;
        RECT 108.300 0.510 108.590 5.800 ;
        RECT 108.930 0.510 109.100 5.380 ;
        RECT 4.270 0.350 5.670 0.510 ;
        RECT 7.510 0.350 11.360 0.510 ;
        RECT 13.020 0.350 16.870 0.510 ;
        RECT 18.660 0.350 20.550 0.510 ;
        RECT 21.980 0.350 23.380 0.510 ;
        RECT 25.220 0.350 29.070 0.510 ;
        RECT 30.730 0.350 34.580 0.510 ;
        RECT 36.370 0.350 38.260 0.510 ;
        RECT 39.690 0.350 41.090 0.510 ;
        RECT 42.930 0.350 46.780 0.510 ;
        RECT 48.440 0.350 52.290 0.510 ;
        RECT 54.080 0.350 55.970 0.510 ;
        RECT 57.400 0.350 58.800 0.510 ;
        RECT 60.640 0.350 64.490 0.510 ;
        RECT 66.150 0.350 70.000 0.510 ;
        RECT 71.790 0.350 73.680 0.510 ;
        RECT 75.110 0.350 76.510 0.510 ;
        RECT 78.350 0.350 82.200 0.510 ;
        RECT 83.860 0.350 87.710 0.510 ;
        RECT 89.500 0.350 91.390 0.510 ;
        RECT 92.820 0.350 94.220 0.510 ;
        RECT 96.060 0.350 99.910 0.510 ;
        RECT 101.570 0.350 105.420 0.510 ;
        RECT 107.210 0.350 109.100 0.510 ;
        RECT 2.680 0.180 109.100 0.350 ;
        RECT 4.270 0.150 5.670 0.180 ;
        RECT 7.510 0.150 11.360 0.180 ;
        RECT 13.020 0.150 16.870 0.180 ;
        RECT 18.660 0.150 20.550 0.180 ;
        RECT 21.980 0.150 23.380 0.180 ;
        RECT 25.220 0.150 29.070 0.180 ;
        RECT 30.730 0.150 34.580 0.180 ;
        RECT 36.370 0.150 38.260 0.180 ;
        RECT 39.690 0.150 41.090 0.180 ;
        RECT 42.930 0.150 46.780 0.180 ;
        RECT 48.440 0.150 52.290 0.180 ;
        RECT 54.080 0.150 55.970 0.180 ;
        RECT 57.400 0.150 58.800 0.180 ;
        RECT 60.640 0.150 64.490 0.180 ;
        RECT 66.150 0.150 70.000 0.180 ;
        RECT 71.790 0.150 73.680 0.180 ;
        RECT 75.110 0.150 76.510 0.180 ;
        RECT 78.350 0.150 82.200 0.180 ;
        RECT 83.860 0.150 87.710 0.180 ;
        RECT 89.500 0.150 91.390 0.180 ;
        RECT 92.820 0.150 94.220 0.180 ;
        RECT 96.060 0.150 99.910 0.180 ;
        RECT 101.570 0.150 105.420 0.180 ;
        RECT 107.210 0.150 109.100 0.180 ;
      LAYER mcon ;
        RECT 11.220 29.360 11.520 29.660 ;
        RECT 11.710 29.360 12.010 29.660 ;
        RECT 12.200 29.360 12.500 29.660 ;
        RECT 12.690 29.360 12.990 29.660 ;
        RECT 14.900 29.360 15.200 29.660 ;
        RECT 15.390 29.360 15.690 29.660 ;
        RECT 15.880 29.360 16.180 29.660 ;
        RECT 16.370 29.360 16.670 29.660 ;
        RECT 16.860 29.360 17.160 29.660 ;
        RECT 17.350 29.360 17.650 29.660 ;
        RECT 17.840 29.360 18.140 29.660 ;
        RECT 18.330 29.360 18.630 29.660 ;
        RECT 20.410 29.360 20.710 29.660 ;
        RECT 20.900 29.360 21.200 29.660 ;
        RECT 21.390 29.360 21.690 29.660 ;
        RECT 21.880 29.360 22.180 29.660 ;
        RECT 22.370 29.360 22.670 29.660 ;
        RECT 22.860 29.360 23.160 29.660 ;
        RECT 23.350 29.360 23.650 29.660 ;
        RECT 23.840 29.360 24.140 29.660 ;
        RECT 26.100 29.360 26.400 29.660 ;
        RECT 26.590 29.360 26.890 29.660 ;
        RECT 27.080 29.360 27.380 29.660 ;
        RECT 28.930 29.360 29.230 29.660 ;
        RECT 29.420 29.360 29.720 29.660 ;
        RECT 29.910 29.360 30.210 29.660 ;
        RECT 30.400 29.360 30.700 29.660 ;
        RECT 32.610 29.360 32.910 29.660 ;
        RECT 33.100 29.360 33.400 29.660 ;
        RECT 33.590 29.360 33.890 29.660 ;
        RECT 34.080 29.360 34.380 29.660 ;
        RECT 34.570 29.360 34.870 29.660 ;
        RECT 35.060 29.360 35.360 29.660 ;
        RECT 35.550 29.360 35.850 29.660 ;
        RECT 36.040 29.360 36.340 29.660 ;
        RECT 38.120 29.360 38.420 29.660 ;
        RECT 38.610 29.360 38.910 29.660 ;
        RECT 39.100 29.360 39.400 29.660 ;
        RECT 39.590 29.360 39.890 29.660 ;
        RECT 40.080 29.360 40.380 29.660 ;
        RECT 40.570 29.360 40.870 29.660 ;
        RECT 41.060 29.360 41.360 29.660 ;
        RECT 41.550 29.360 41.850 29.660 ;
        RECT 43.810 29.360 44.110 29.660 ;
        RECT 44.300 29.360 44.600 29.660 ;
        RECT 44.790 29.360 45.090 29.660 ;
        RECT 46.640 29.360 46.940 29.660 ;
        RECT 47.130 29.360 47.430 29.660 ;
        RECT 47.620 29.360 47.920 29.660 ;
        RECT 48.110 29.360 48.410 29.660 ;
        RECT 50.320 29.360 50.620 29.660 ;
        RECT 50.810 29.360 51.110 29.660 ;
        RECT 51.300 29.360 51.600 29.660 ;
        RECT 51.790 29.360 52.090 29.660 ;
        RECT 52.280 29.360 52.580 29.660 ;
        RECT 52.770 29.360 53.070 29.660 ;
        RECT 53.260 29.360 53.560 29.660 ;
        RECT 53.750 29.360 54.050 29.660 ;
        RECT 55.830 29.360 56.130 29.660 ;
        RECT 56.320 29.360 56.620 29.660 ;
        RECT 56.810 29.360 57.110 29.660 ;
        RECT 57.300 29.360 57.600 29.660 ;
        RECT 57.790 29.360 58.090 29.660 ;
        RECT 58.280 29.360 58.580 29.660 ;
        RECT 58.770 29.360 59.070 29.660 ;
        RECT 59.260 29.360 59.560 29.660 ;
        RECT 61.520 29.360 61.820 29.660 ;
        RECT 62.010 29.360 62.310 29.660 ;
        RECT 62.500 29.360 62.800 29.660 ;
        RECT 64.350 29.360 64.650 29.660 ;
        RECT 64.840 29.360 65.140 29.660 ;
        RECT 65.330 29.360 65.630 29.660 ;
        RECT 65.820 29.360 66.120 29.660 ;
        RECT 68.030 29.360 68.330 29.660 ;
        RECT 68.520 29.360 68.820 29.660 ;
        RECT 69.010 29.360 69.310 29.660 ;
        RECT 69.500 29.360 69.800 29.660 ;
        RECT 69.990 29.360 70.290 29.660 ;
        RECT 70.480 29.360 70.780 29.660 ;
        RECT 70.970 29.360 71.270 29.660 ;
        RECT 71.460 29.360 71.760 29.660 ;
        RECT 73.540 29.360 73.840 29.660 ;
        RECT 74.030 29.360 74.330 29.660 ;
        RECT 74.520 29.360 74.820 29.660 ;
        RECT 75.010 29.360 75.310 29.660 ;
        RECT 75.500 29.360 75.800 29.660 ;
        RECT 75.990 29.360 76.290 29.660 ;
        RECT 76.480 29.360 76.780 29.660 ;
        RECT 76.970 29.360 77.270 29.660 ;
        RECT 79.230 29.360 79.530 29.660 ;
        RECT 79.720 29.360 80.020 29.660 ;
        RECT 80.210 29.360 80.510 29.660 ;
        RECT 82.060 29.360 82.360 29.660 ;
        RECT 82.550 29.360 82.850 29.660 ;
        RECT 83.040 29.360 83.340 29.660 ;
        RECT 83.530 29.360 83.830 29.660 ;
        RECT 85.740 29.360 86.040 29.660 ;
        RECT 86.230 29.360 86.530 29.660 ;
        RECT 86.720 29.360 87.020 29.660 ;
        RECT 87.210 29.360 87.510 29.660 ;
        RECT 87.700 29.360 88.000 29.660 ;
        RECT 88.190 29.360 88.490 29.660 ;
        RECT 88.680 29.360 88.980 29.660 ;
        RECT 89.170 29.360 89.470 29.660 ;
        RECT 91.250 29.360 91.550 29.660 ;
        RECT 91.740 29.360 92.040 29.660 ;
        RECT 92.230 29.360 92.530 29.660 ;
        RECT 92.720 29.360 93.020 29.660 ;
        RECT 93.210 29.360 93.510 29.660 ;
        RECT 93.700 29.360 94.000 29.660 ;
        RECT 94.190 29.360 94.490 29.660 ;
        RECT 94.680 29.360 94.980 29.660 ;
        RECT 96.940 29.360 97.240 29.660 ;
        RECT 97.430 29.360 97.730 29.660 ;
        RECT 97.920 29.360 98.220 29.660 ;
        RECT 1.835 25.435 2.005 25.605 ;
        RECT 2.295 25.435 2.465 25.605 ;
        RECT 2.755 25.435 2.925 25.605 ;
        RECT 3.215 25.435 3.385 25.605 ;
        RECT 3.675 25.435 3.845 25.605 ;
        RECT 5.830 25.435 6.000 25.605 ;
        RECT 6.290 25.435 6.460 25.605 ;
        RECT 6.750 25.435 6.920 25.605 ;
        RECT 4.330 0.180 4.630 0.480 ;
        RECT 4.820 0.180 5.120 0.480 ;
        RECT 5.310 0.180 5.610 0.480 ;
        RECT 7.570 0.180 7.870 0.480 ;
        RECT 8.060 0.180 8.360 0.480 ;
        RECT 8.550 0.180 8.850 0.480 ;
        RECT 9.040 0.180 9.340 0.480 ;
        RECT 9.530 0.180 9.830 0.480 ;
        RECT 10.020 0.180 10.320 0.480 ;
        RECT 10.510 0.180 10.810 0.480 ;
        RECT 11.000 0.180 11.300 0.480 ;
        RECT 13.080 0.180 13.380 0.480 ;
        RECT 13.570 0.180 13.870 0.480 ;
        RECT 14.060 0.180 14.360 0.480 ;
        RECT 14.550 0.180 14.850 0.480 ;
        RECT 15.040 0.180 15.340 0.480 ;
        RECT 15.530 0.180 15.830 0.480 ;
        RECT 16.020 0.180 16.320 0.480 ;
        RECT 16.510 0.180 16.810 0.480 ;
        RECT 18.720 0.180 19.020 0.480 ;
        RECT 19.210 0.180 19.510 0.480 ;
        RECT 19.700 0.180 20.000 0.480 ;
        RECT 20.190 0.180 20.490 0.480 ;
        RECT 22.040 0.180 22.340 0.480 ;
        RECT 22.530 0.180 22.830 0.480 ;
        RECT 23.020 0.180 23.320 0.480 ;
        RECT 25.280 0.180 25.580 0.480 ;
        RECT 25.770 0.180 26.070 0.480 ;
        RECT 26.260 0.180 26.560 0.480 ;
        RECT 26.750 0.180 27.050 0.480 ;
        RECT 27.240 0.180 27.540 0.480 ;
        RECT 27.730 0.180 28.030 0.480 ;
        RECT 28.220 0.180 28.520 0.480 ;
        RECT 28.710 0.180 29.010 0.480 ;
        RECT 30.790 0.180 31.090 0.480 ;
        RECT 31.280 0.180 31.580 0.480 ;
        RECT 31.770 0.180 32.070 0.480 ;
        RECT 32.260 0.180 32.560 0.480 ;
        RECT 32.750 0.180 33.050 0.480 ;
        RECT 33.240 0.180 33.540 0.480 ;
        RECT 33.730 0.180 34.030 0.480 ;
        RECT 34.220 0.180 34.520 0.480 ;
        RECT 36.430 0.180 36.730 0.480 ;
        RECT 36.920 0.180 37.220 0.480 ;
        RECT 37.410 0.180 37.710 0.480 ;
        RECT 37.900 0.180 38.200 0.480 ;
        RECT 39.750 0.180 40.050 0.480 ;
        RECT 40.240 0.180 40.540 0.480 ;
        RECT 40.730 0.180 41.030 0.480 ;
        RECT 42.990 0.180 43.290 0.480 ;
        RECT 43.480 0.180 43.780 0.480 ;
        RECT 43.970 0.180 44.270 0.480 ;
        RECT 44.460 0.180 44.760 0.480 ;
        RECT 44.950 0.180 45.250 0.480 ;
        RECT 45.440 0.180 45.740 0.480 ;
        RECT 45.930 0.180 46.230 0.480 ;
        RECT 46.420 0.180 46.720 0.480 ;
        RECT 48.500 0.180 48.800 0.480 ;
        RECT 48.990 0.180 49.290 0.480 ;
        RECT 49.480 0.180 49.780 0.480 ;
        RECT 49.970 0.180 50.270 0.480 ;
        RECT 50.460 0.180 50.760 0.480 ;
        RECT 50.950 0.180 51.250 0.480 ;
        RECT 51.440 0.180 51.740 0.480 ;
        RECT 51.930 0.180 52.230 0.480 ;
        RECT 54.140 0.180 54.440 0.480 ;
        RECT 54.630 0.180 54.930 0.480 ;
        RECT 55.120 0.180 55.420 0.480 ;
        RECT 55.610 0.180 55.910 0.480 ;
        RECT 57.460 0.180 57.760 0.480 ;
        RECT 57.950 0.180 58.250 0.480 ;
        RECT 58.440 0.180 58.740 0.480 ;
        RECT 60.700 0.180 61.000 0.480 ;
        RECT 61.190 0.180 61.490 0.480 ;
        RECT 61.680 0.180 61.980 0.480 ;
        RECT 62.170 0.180 62.470 0.480 ;
        RECT 62.660 0.180 62.960 0.480 ;
        RECT 63.150 0.180 63.450 0.480 ;
        RECT 63.640 0.180 63.940 0.480 ;
        RECT 64.130 0.180 64.430 0.480 ;
        RECT 66.210 0.180 66.510 0.480 ;
        RECT 66.700 0.180 67.000 0.480 ;
        RECT 67.190 0.180 67.490 0.480 ;
        RECT 67.680 0.180 67.980 0.480 ;
        RECT 68.170 0.180 68.470 0.480 ;
        RECT 68.660 0.180 68.960 0.480 ;
        RECT 69.150 0.180 69.450 0.480 ;
        RECT 69.640 0.180 69.940 0.480 ;
        RECT 71.850 0.180 72.150 0.480 ;
        RECT 72.340 0.180 72.640 0.480 ;
        RECT 72.830 0.180 73.130 0.480 ;
        RECT 73.320 0.180 73.620 0.480 ;
        RECT 75.170 0.180 75.470 0.480 ;
        RECT 75.660 0.180 75.960 0.480 ;
        RECT 76.150 0.180 76.450 0.480 ;
        RECT 78.410 0.180 78.710 0.480 ;
        RECT 78.900 0.180 79.200 0.480 ;
        RECT 79.390 0.180 79.690 0.480 ;
        RECT 79.880 0.180 80.180 0.480 ;
        RECT 80.370 0.180 80.670 0.480 ;
        RECT 80.860 0.180 81.160 0.480 ;
        RECT 81.350 0.180 81.650 0.480 ;
        RECT 81.840 0.180 82.140 0.480 ;
        RECT 83.920 0.180 84.220 0.480 ;
        RECT 84.410 0.180 84.710 0.480 ;
        RECT 84.900 0.180 85.200 0.480 ;
        RECT 85.390 0.180 85.690 0.480 ;
        RECT 85.880 0.180 86.180 0.480 ;
        RECT 86.370 0.180 86.670 0.480 ;
        RECT 86.860 0.180 87.160 0.480 ;
        RECT 87.350 0.180 87.650 0.480 ;
        RECT 89.560 0.180 89.860 0.480 ;
        RECT 90.050 0.180 90.350 0.480 ;
        RECT 90.540 0.180 90.840 0.480 ;
        RECT 91.030 0.180 91.330 0.480 ;
        RECT 92.880 0.180 93.180 0.480 ;
        RECT 93.370 0.180 93.670 0.480 ;
        RECT 93.860 0.180 94.160 0.480 ;
        RECT 96.120 0.180 96.420 0.480 ;
        RECT 96.610 0.180 96.910 0.480 ;
        RECT 97.100 0.180 97.400 0.480 ;
        RECT 97.590 0.180 97.890 0.480 ;
        RECT 98.080 0.180 98.380 0.480 ;
        RECT 98.570 0.180 98.870 0.480 ;
        RECT 99.060 0.180 99.360 0.480 ;
        RECT 99.550 0.180 99.850 0.480 ;
        RECT 101.630 0.180 101.930 0.480 ;
        RECT 102.120 0.180 102.420 0.480 ;
        RECT 102.610 0.180 102.910 0.480 ;
        RECT 103.100 0.180 103.400 0.480 ;
        RECT 103.590 0.180 103.890 0.480 ;
        RECT 104.080 0.180 104.380 0.480 ;
        RECT 104.570 0.180 104.870 0.480 ;
        RECT 105.060 0.180 105.360 0.480 ;
        RECT 107.270 0.180 107.570 0.480 ;
        RECT 107.760 0.180 108.060 0.480 ;
        RECT 108.250 0.180 108.550 0.480 ;
        RECT 108.740 0.180 109.040 0.480 ;
      LAYER met1 ;
        RECT 10.900 29.270 100.050 29.750 ;
        RECT -5.000 25.280 7.065 25.760 ;
        RECT 2.500 0.090 109.280 0.570 ;
      LAYER via ;
        RECT 13.130 29.360 13.430 29.660 ;
        RECT 13.490 29.360 13.790 29.660 ;
        RECT 13.850 29.360 14.150 29.660 ;
        RECT 14.210 29.360 14.510 29.660 ;
        RECT 14.570 29.360 14.870 29.660 ;
        RECT 41.130 29.360 41.430 29.660 ;
        RECT 41.490 29.360 41.790 29.660 ;
        RECT 41.850 29.360 42.150 29.660 ;
        RECT 42.210 29.360 42.510 29.660 ;
        RECT 42.570 29.360 42.870 29.660 ;
        RECT 69.130 29.360 69.430 29.660 ;
        RECT 69.490 29.360 69.790 29.660 ;
        RECT 69.850 29.360 70.150 29.660 ;
        RECT 70.210 29.360 70.510 29.660 ;
        RECT 70.570 29.360 70.870 29.660 ;
        RECT 97.130 29.360 97.430 29.660 ;
        RECT 97.490 29.360 97.790 29.660 ;
        RECT 97.850 29.360 98.150 29.660 ;
        RECT 98.210 29.360 98.510 29.660 ;
        RECT 98.570 29.360 98.870 29.660 ;
        RECT -4.870 25.370 -4.570 25.670 ;
        RECT -4.510 25.370 -4.210 25.670 ;
        RECT -4.150 25.370 -3.850 25.670 ;
        RECT -3.790 25.370 -3.490 25.670 ;
        RECT -3.430 25.370 -3.130 25.670 ;
        RECT 13.130 0.180 13.430 0.480 ;
        RECT 13.490 0.180 13.790 0.480 ;
        RECT 13.850 0.180 14.150 0.480 ;
        RECT 14.210 0.180 14.510 0.480 ;
        RECT 14.570 0.180 14.870 0.480 ;
        RECT 41.130 0.180 41.430 0.480 ;
        RECT 41.490 0.180 41.790 0.480 ;
        RECT 41.850 0.180 42.150 0.480 ;
        RECT 42.210 0.180 42.510 0.480 ;
        RECT 42.570 0.180 42.870 0.480 ;
        RECT 69.130 0.180 69.430 0.480 ;
        RECT 69.490 0.180 69.790 0.480 ;
        RECT 69.850 0.180 70.150 0.480 ;
        RECT 70.210 0.180 70.510 0.480 ;
        RECT 70.570 0.180 70.870 0.480 ;
        RECT 97.130 0.180 97.430 0.480 ;
        RECT 97.490 0.180 97.790 0.480 ;
        RECT 97.850 0.180 98.150 0.480 ;
        RECT 98.210 0.180 98.510 0.480 ;
        RECT 98.570 0.180 98.870 0.480 ;
      LAYER met2 ;
        RECT 13.000 29.270 15.000 29.750 ;
        RECT 41.000 29.270 43.000 29.750 ;
        RECT 69.000 29.270 71.000 29.750 ;
        RECT 97.000 29.270 99.000 29.750 ;
        RECT -5.000 25.280 -3.000 25.760 ;
        RECT 13.000 0.090 15.000 0.570 ;
        RECT 41.000 0.090 43.000 0.570 ;
        RECT 69.000 0.090 71.000 0.570 ;
        RECT 97.000 0.090 99.000 0.570 ;
      LAYER via2 ;
        RECT 13.180 29.350 13.500 29.670 ;
        RECT 13.620 29.350 13.940 29.670 ;
        RECT 14.060 29.350 14.380 29.670 ;
        RECT 14.500 29.350 14.820 29.670 ;
        RECT 41.180 29.350 41.500 29.670 ;
        RECT 41.620 29.350 41.940 29.670 ;
        RECT 42.060 29.350 42.380 29.670 ;
        RECT 42.500 29.350 42.820 29.670 ;
        RECT 69.180 29.350 69.500 29.670 ;
        RECT 69.620 29.350 69.940 29.670 ;
        RECT 70.060 29.350 70.380 29.670 ;
        RECT 70.500 29.350 70.820 29.670 ;
        RECT 97.180 29.350 97.500 29.670 ;
        RECT 97.620 29.350 97.940 29.670 ;
        RECT 98.060 29.350 98.380 29.670 ;
        RECT 98.500 29.350 98.820 29.670 ;
        RECT -4.820 25.360 -4.500 25.680 ;
        RECT -4.380 25.360 -4.060 25.680 ;
        RECT -3.940 25.360 -3.620 25.680 ;
        RECT -3.500 25.360 -3.180 25.680 ;
        RECT 13.180 0.170 13.500 0.490 ;
        RECT 13.620 0.170 13.940 0.490 ;
        RECT 14.060 0.170 14.380 0.490 ;
        RECT 14.500 0.170 14.820 0.490 ;
        RECT 41.180 0.170 41.500 0.490 ;
        RECT 41.620 0.170 41.940 0.490 ;
        RECT 42.060 0.170 42.380 0.490 ;
        RECT 42.500 0.170 42.820 0.490 ;
        RECT 69.180 0.170 69.500 0.490 ;
        RECT 69.620 0.170 69.940 0.490 ;
        RECT 70.060 0.170 70.380 0.490 ;
        RECT 70.500 0.170 70.820 0.490 ;
        RECT 97.180 0.170 97.500 0.490 ;
        RECT 97.620 0.170 97.940 0.490 ;
        RECT 98.060 0.170 98.380 0.490 ;
        RECT 98.500 0.170 98.820 0.490 ;
      LAYER met3 ;
        RECT -5.000 65.000 117.000 67.000 ;
        RECT 13.000 29.270 15.000 29.750 ;
        RECT 41.000 29.270 43.000 29.750 ;
        RECT 69.000 29.270 71.000 29.750 ;
        RECT 97.000 29.270 99.000 29.750 ;
        RECT -5.000 25.280 -3.000 25.760 ;
        RECT 13.000 0.090 15.000 0.570 ;
        RECT 41.000 0.090 43.000 0.570 ;
        RECT 69.000 0.090 71.000 0.570 ;
        RECT 97.000 0.090 99.000 0.570 ;
        RECT -5.000 -38.000 117.000 -36.000 ;
      LAYER via3 ;
        RECT -4.800 66.400 -4.400 66.800 ;
        RECT -4.200 66.400 -3.800 66.800 ;
        RECT -3.600 66.400 -3.200 66.800 ;
        RECT 13.200 66.400 13.600 66.800 ;
        RECT 13.800 66.400 14.200 66.800 ;
        RECT 14.400 66.400 14.800 66.800 ;
        RECT 41.200 66.400 41.600 66.800 ;
        RECT 41.800 66.400 42.200 66.800 ;
        RECT 42.400 66.400 42.800 66.800 ;
        RECT 69.200 66.400 69.600 66.800 ;
        RECT 69.800 66.400 70.200 66.800 ;
        RECT 70.400 66.400 70.800 66.800 ;
        RECT 97.200 66.400 97.600 66.800 ;
        RECT 97.800 66.400 98.200 66.800 ;
        RECT 98.400 66.400 98.800 66.800 ;
        RECT 115.200 66.400 115.600 66.800 ;
        RECT 115.800 66.400 116.200 66.800 ;
        RECT 116.400 66.400 116.800 66.800 ;
        RECT -4.800 65.800 -4.400 66.200 ;
        RECT -4.200 65.800 -3.800 66.200 ;
        RECT -3.600 65.800 -3.200 66.200 ;
        RECT 13.200 65.800 13.600 66.200 ;
        RECT 13.800 65.800 14.200 66.200 ;
        RECT 14.400 65.800 14.800 66.200 ;
        RECT 41.200 65.800 41.600 66.200 ;
        RECT 41.800 65.800 42.200 66.200 ;
        RECT 42.400 65.800 42.800 66.200 ;
        RECT 69.200 65.800 69.600 66.200 ;
        RECT 69.800 65.800 70.200 66.200 ;
        RECT 70.400 65.800 70.800 66.200 ;
        RECT 97.200 65.800 97.600 66.200 ;
        RECT 97.800 65.800 98.200 66.200 ;
        RECT 98.400 65.800 98.800 66.200 ;
        RECT 115.200 65.800 115.600 66.200 ;
        RECT 115.800 65.800 116.200 66.200 ;
        RECT 116.400 65.800 116.800 66.200 ;
        RECT -4.800 65.200 -4.400 65.600 ;
        RECT -4.200 65.200 -3.800 65.600 ;
        RECT -3.600 65.200 -3.200 65.600 ;
        RECT 13.200 65.200 13.600 65.600 ;
        RECT 13.800 65.200 14.200 65.600 ;
        RECT 14.400 65.200 14.800 65.600 ;
        RECT 41.200 65.200 41.600 65.600 ;
        RECT 41.800 65.200 42.200 65.600 ;
        RECT 42.400 65.200 42.800 65.600 ;
        RECT 69.200 65.200 69.600 65.600 ;
        RECT 69.800 65.200 70.200 65.600 ;
        RECT 70.400 65.200 70.800 65.600 ;
        RECT 97.200 65.200 97.600 65.600 ;
        RECT 97.800 65.200 98.200 65.600 ;
        RECT 98.400 65.200 98.800 65.600 ;
        RECT 115.200 65.200 115.600 65.600 ;
        RECT 115.800 65.200 116.200 65.600 ;
        RECT 116.400 65.200 116.800 65.600 ;
        RECT 13.160 29.330 13.520 29.695 ;
        RECT 13.600 29.330 13.960 29.695 ;
        RECT 14.040 29.330 14.400 29.695 ;
        RECT 14.480 29.330 14.840 29.695 ;
        RECT 41.160 29.330 41.520 29.695 ;
        RECT 41.600 29.330 41.960 29.695 ;
        RECT 42.040 29.330 42.400 29.695 ;
        RECT 42.480 29.330 42.840 29.695 ;
        RECT 69.160 29.330 69.520 29.695 ;
        RECT 69.600 29.330 69.960 29.695 ;
        RECT 70.040 29.330 70.400 29.695 ;
        RECT 70.480 29.330 70.840 29.695 ;
        RECT 97.160 29.330 97.520 29.695 ;
        RECT 97.600 29.330 97.960 29.695 ;
        RECT 98.040 29.330 98.400 29.695 ;
        RECT 98.480 29.330 98.840 29.695 ;
        RECT -4.840 25.340 -4.480 25.705 ;
        RECT -4.400 25.340 -4.040 25.705 ;
        RECT -3.960 25.340 -3.600 25.705 ;
        RECT -3.520 25.340 -3.160 25.705 ;
        RECT 13.160 0.150 13.520 0.515 ;
        RECT 13.600 0.150 13.960 0.515 ;
        RECT 14.040 0.150 14.400 0.515 ;
        RECT 14.480 0.150 14.840 0.515 ;
        RECT 41.160 0.150 41.520 0.515 ;
        RECT 41.600 0.150 41.960 0.515 ;
        RECT 42.040 0.150 42.400 0.515 ;
        RECT 42.480 0.150 42.840 0.515 ;
        RECT 69.160 0.150 69.520 0.515 ;
        RECT 69.600 0.150 69.960 0.515 ;
        RECT 70.040 0.150 70.400 0.515 ;
        RECT 70.480 0.150 70.840 0.515 ;
        RECT 97.160 0.150 97.520 0.515 ;
        RECT 97.600 0.150 97.960 0.515 ;
        RECT 98.040 0.150 98.400 0.515 ;
        RECT 98.480 0.150 98.840 0.515 ;
        RECT -4.800 -36.600 -4.400 -36.200 ;
        RECT -4.200 -36.600 -3.800 -36.200 ;
        RECT -3.600 -36.600 -3.200 -36.200 ;
        RECT 13.200 -36.600 13.600 -36.200 ;
        RECT 13.800 -36.600 14.200 -36.200 ;
        RECT 14.400 -36.600 14.800 -36.200 ;
        RECT 41.200 -36.600 41.600 -36.200 ;
        RECT 41.800 -36.600 42.200 -36.200 ;
        RECT 42.400 -36.600 42.800 -36.200 ;
        RECT 69.200 -36.600 69.600 -36.200 ;
        RECT 69.800 -36.600 70.200 -36.200 ;
        RECT 70.400 -36.600 70.800 -36.200 ;
        RECT 97.200 -36.600 97.600 -36.200 ;
        RECT 97.800 -36.600 98.200 -36.200 ;
        RECT 98.400 -36.600 98.800 -36.200 ;
        RECT 115.200 -36.600 115.600 -36.200 ;
        RECT 115.800 -36.600 116.200 -36.200 ;
        RECT 116.400 -36.600 116.800 -36.200 ;
        RECT -4.800 -37.200 -4.400 -36.800 ;
        RECT -4.200 -37.200 -3.800 -36.800 ;
        RECT -3.600 -37.200 -3.200 -36.800 ;
        RECT 13.200 -37.200 13.600 -36.800 ;
        RECT 13.800 -37.200 14.200 -36.800 ;
        RECT 14.400 -37.200 14.800 -36.800 ;
        RECT 41.200 -37.200 41.600 -36.800 ;
        RECT 41.800 -37.200 42.200 -36.800 ;
        RECT 42.400 -37.200 42.800 -36.800 ;
        RECT 69.200 -37.200 69.600 -36.800 ;
        RECT 69.800 -37.200 70.200 -36.800 ;
        RECT 70.400 -37.200 70.800 -36.800 ;
        RECT 97.200 -37.200 97.600 -36.800 ;
        RECT 97.800 -37.200 98.200 -36.800 ;
        RECT 98.400 -37.200 98.800 -36.800 ;
        RECT 115.200 -37.200 115.600 -36.800 ;
        RECT 115.800 -37.200 116.200 -36.800 ;
        RECT 116.400 -37.200 116.800 -36.800 ;
        RECT -4.800 -37.800 -4.400 -37.400 ;
        RECT -4.200 -37.800 -3.800 -37.400 ;
        RECT -3.600 -37.800 -3.200 -37.400 ;
        RECT 13.200 -37.800 13.600 -37.400 ;
        RECT 13.800 -37.800 14.200 -37.400 ;
        RECT 14.400 -37.800 14.800 -37.400 ;
        RECT 41.200 -37.800 41.600 -37.400 ;
        RECT 41.800 -37.800 42.200 -37.400 ;
        RECT 42.400 -37.800 42.800 -37.400 ;
        RECT 69.200 -37.800 69.600 -37.400 ;
        RECT 69.800 -37.800 70.200 -37.400 ;
        RECT 70.400 -37.800 70.800 -37.400 ;
        RECT 97.200 -37.800 97.600 -37.400 ;
        RECT 97.800 -37.800 98.200 -37.400 ;
        RECT 98.400 -37.800 98.800 -37.400 ;
        RECT 115.200 -37.800 115.600 -37.400 ;
        RECT 115.800 -37.800 116.200 -37.400 ;
        RECT 116.400 -37.800 116.800 -37.400 ;
      LAYER met4 ;
        RECT -5.000 -38.000 -3.000 67.000 ;
        RECT 13.000 -38.000 15.000 67.000 ;
        RECT 41.000 -38.000 43.000 67.000 ;
        RECT 69.000 -38.000 71.000 67.000 ;
        RECT 97.000 -38.000 99.000 67.000 ;
        RECT 115.000 -38.000 117.000 67.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 10.000 30.700 101.000 31.000 ;
        RECT 2.205 22.885 3.140 23.285 ;
        RECT 6.460 22.885 6.800 23.545 ;
        RECT 1.690 22.715 3.990 22.885 ;
        RECT 5.685 22.715 7.065 22.885 ;
        RECT 10.000 15.070 10.300 30.700 ;
        RECT 100.700 15.070 101.000 30.700 ;
        RECT 103.500 24.015 105.500 24.380 ;
        RECT 1.700 14.770 110.825 15.070 ;
        RECT 1.700 -0.800 2.000 14.770 ;
        RECT 110.500 14.700 110.825 14.770 ;
        RECT 110.500 -0.800 110.800 14.700 ;
        RECT 1.700 -1.100 110.800 -0.800 ;
      LAYER mcon ;
        RECT 27.110 30.700 27.410 31.000 ;
        RECT 27.600 30.700 27.900 31.000 ;
        RECT 28.100 30.700 28.400 31.000 ;
        RECT 28.590 30.700 28.890 31.000 ;
        RECT 55.110 30.700 55.410 31.000 ;
        RECT 55.600 30.700 55.900 31.000 ;
        RECT 56.100 30.700 56.400 31.000 ;
        RECT 56.590 30.700 56.890 31.000 ;
        RECT 83.110 30.700 83.410 31.000 ;
        RECT 83.600 30.700 83.900 31.000 ;
        RECT 84.100 30.700 84.400 31.000 ;
        RECT 84.590 30.700 84.890 31.000 ;
        RECT 1.835 22.715 2.005 22.885 ;
        RECT 2.295 22.715 2.465 22.885 ;
        RECT 2.755 22.715 2.925 22.885 ;
        RECT 3.215 22.715 3.385 22.885 ;
        RECT 3.675 22.715 3.845 22.885 ;
        RECT 5.830 22.715 6.000 22.885 ;
        RECT 6.290 22.715 6.460 22.885 ;
        RECT 6.750 22.715 6.920 22.885 ;
        RECT 103.600 24.050 103.900 24.350 ;
        RECT 104.100 24.050 104.400 24.350 ;
        RECT 104.600 24.050 104.900 24.350 ;
        RECT 105.100 24.050 105.400 24.350 ;
        RECT 27.110 -1.100 27.410 -0.800 ;
        RECT 27.600 -1.100 27.900 -0.800 ;
        RECT 28.100 -1.100 28.400 -0.800 ;
        RECT 28.590 -1.100 28.890 -0.800 ;
        RECT 55.110 -1.100 55.410 -0.800 ;
        RECT 55.600 -1.100 55.900 -0.800 ;
        RECT 56.100 -1.100 56.400 -0.800 ;
        RECT 56.590 -1.100 56.890 -0.800 ;
      LAYER met1 ;
        RECT 27.080 30.610 28.920 31.090 ;
        RECT 55.080 30.610 56.920 31.090 ;
        RECT 83.080 30.610 84.920 31.090 ;
        RECT 111.130 24.380 112.870 24.440 ;
        RECT 103.500 24.020 113.000 24.380 ;
        RECT 103.500 24.015 105.505 24.020 ;
        RECT 111.130 23.960 112.870 24.020 ;
        RECT -1.000 22.560 7.065 23.040 ;
        RECT 27.080 -1.190 28.920 -0.710 ;
        RECT 55.080 -1.190 56.920 -0.710 ;
      LAYER via ;
        RECT 27.130 30.700 27.430 31.000 ;
        RECT 27.490 30.700 27.790 31.000 ;
        RECT 27.850 30.700 28.150 31.000 ;
        RECT 28.210 30.700 28.510 31.000 ;
        RECT 28.570 30.700 28.870 31.000 ;
        RECT 55.130 30.700 55.430 31.000 ;
        RECT 55.490 30.700 55.790 31.000 ;
        RECT 55.850 30.700 56.150 31.000 ;
        RECT 56.210 30.700 56.510 31.000 ;
        RECT 56.570 30.700 56.870 31.000 ;
        RECT 83.130 30.700 83.430 31.000 ;
        RECT 83.490 30.700 83.790 31.000 ;
        RECT 83.850 30.700 84.150 31.000 ;
        RECT 84.210 30.700 84.510 31.000 ;
        RECT 84.570 30.700 84.870 31.000 ;
        RECT 111.130 24.050 111.430 24.350 ;
        RECT 111.490 24.050 111.790 24.350 ;
        RECT 111.850 24.050 112.150 24.350 ;
        RECT 112.210 24.050 112.510 24.350 ;
        RECT 112.570 24.050 112.870 24.350 ;
        RECT -0.870 22.650 -0.570 22.950 ;
        RECT -0.510 22.650 -0.210 22.950 ;
        RECT -0.150 22.650 0.150 22.950 ;
        RECT 0.210 22.650 0.510 22.950 ;
        RECT 0.570 22.650 0.870 22.950 ;
        RECT 27.130 -1.100 27.430 -0.800 ;
        RECT 27.490 -1.100 27.790 -0.800 ;
        RECT 27.850 -1.100 28.150 -0.800 ;
        RECT 28.210 -1.100 28.510 -0.800 ;
        RECT 28.570 -1.100 28.870 -0.800 ;
        RECT 55.130 -1.100 55.430 -0.800 ;
        RECT 55.490 -1.100 55.790 -0.800 ;
        RECT 55.850 -1.100 56.150 -0.800 ;
        RECT 56.210 -1.100 56.510 -0.800 ;
        RECT 56.570 -1.100 56.870 -0.800 ;
      LAYER met2 ;
        RECT 27.000 30.610 29.000 31.090 ;
        RECT 55.000 30.610 57.000 31.090 ;
        RECT 83.000 30.610 85.000 31.090 ;
        RECT 111.000 23.960 113.000 24.440 ;
        RECT -1.000 22.560 1.000 23.040 ;
        RECT 27.000 -1.190 29.000 -0.710 ;
        RECT 55.000 -1.190 57.000 -0.710 ;
      LAYER via2 ;
        RECT 27.180 30.690 27.500 31.010 ;
        RECT 27.620 30.690 27.940 31.010 ;
        RECT 28.060 30.690 28.380 31.010 ;
        RECT 28.500 30.690 28.820 31.010 ;
        RECT 55.180 30.690 55.500 31.010 ;
        RECT 55.620 30.690 55.940 31.010 ;
        RECT 56.060 30.690 56.380 31.010 ;
        RECT 56.500 30.690 56.820 31.010 ;
        RECT 83.180 30.690 83.500 31.010 ;
        RECT 83.620 30.690 83.940 31.010 ;
        RECT 84.060 30.690 84.380 31.010 ;
        RECT 84.500 30.690 84.820 31.010 ;
        RECT 111.180 24.040 111.500 24.360 ;
        RECT 111.620 24.040 111.940 24.360 ;
        RECT 112.060 24.040 112.380 24.360 ;
        RECT 112.500 24.040 112.820 24.360 ;
        RECT -0.820 22.640 -0.500 22.960 ;
        RECT -0.380 22.640 -0.060 22.960 ;
        RECT 0.060 22.640 0.380 22.960 ;
        RECT 0.500 22.640 0.820 22.960 ;
        RECT 27.180 -1.110 27.500 -0.790 ;
        RECT 27.620 -1.110 27.940 -0.790 ;
        RECT 28.060 -1.110 28.380 -0.790 ;
        RECT 28.500 -1.110 28.820 -0.790 ;
        RECT 55.180 -1.110 55.500 -0.790 ;
        RECT 55.620 -1.110 55.940 -0.790 ;
        RECT 56.060 -1.110 56.380 -0.790 ;
        RECT 56.500 -1.110 56.820 -0.790 ;
      LAYER met3 ;
        RECT -1.000 61.000 113.000 63.000 ;
        RECT 27.000 30.610 29.000 31.090 ;
        RECT 55.000 30.610 57.000 31.090 ;
        RECT 83.000 30.610 85.000 31.090 ;
        RECT 111.000 23.960 113.000 24.440 ;
        RECT -1.000 22.560 1.000 23.040 ;
        RECT 27.000 -1.190 29.000 -0.710 ;
        RECT 55.000 -1.190 57.000 -0.710 ;
        RECT -1.000 -34.000 113.000 -32.000 ;
      LAYER via3 ;
        RECT -0.800 62.400 -0.400 62.800 ;
        RECT -0.200 62.400 0.200 62.800 ;
        RECT 0.400 62.400 0.800 62.800 ;
        RECT 27.200 62.400 27.600 62.800 ;
        RECT 27.800 62.400 28.200 62.800 ;
        RECT 28.400 62.400 28.800 62.800 ;
        RECT 55.200 62.400 55.600 62.800 ;
        RECT 55.800 62.400 56.200 62.800 ;
        RECT 56.400 62.400 56.800 62.800 ;
        RECT 83.200 62.400 83.600 62.800 ;
        RECT 83.800 62.400 84.200 62.800 ;
        RECT 84.400 62.400 84.800 62.800 ;
        RECT 111.200 62.400 111.600 62.800 ;
        RECT 111.800 62.400 112.200 62.800 ;
        RECT 112.400 62.400 112.800 62.800 ;
        RECT -0.800 61.800 -0.400 62.200 ;
        RECT -0.200 61.800 0.200 62.200 ;
        RECT 0.400 61.800 0.800 62.200 ;
        RECT 27.200 61.800 27.600 62.200 ;
        RECT 27.800 61.800 28.200 62.200 ;
        RECT 28.400 61.800 28.800 62.200 ;
        RECT 55.200 61.800 55.600 62.200 ;
        RECT 55.800 61.800 56.200 62.200 ;
        RECT 56.400 61.800 56.800 62.200 ;
        RECT 83.200 61.800 83.600 62.200 ;
        RECT 83.800 61.800 84.200 62.200 ;
        RECT 84.400 61.800 84.800 62.200 ;
        RECT 111.200 61.800 111.600 62.200 ;
        RECT 111.800 61.800 112.200 62.200 ;
        RECT 112.400 61.800 112.800 62.200 ;
        RECT -0.800 61.200 -0.400 61.600 ;
        RECT -0.200 61.200 0.200 61.600 ;
        RECT 0.400 61.200 0.800 61.600 ;
        RECT 27.200 61.200 27.600 61.600 ;
        RECT 27.800 61.200 28.200 61.600 ;
        RECT 28.400 61.200 28.800 61.600 ;
        RECT 55.200 61.200 55.600 61.600 ;
        RECT 55.800 61.200 56.200 61.600 ;
        RECT 56.400 61.200 56.800 61.600 ;
        RECT 83.200 61.200 83.600 61.600 ;
        RECT 83.800 61.200 84.200 61.600 ;
        RECT 84.400 61.200 84.800 61.600 ;
        RECT 111.200 61.200 111.600 61.600 ;
        RECT 111.800 61.200 112.200 61.600 ;
        RECT 112.400 61.200 112.800 61.600 ;
        RECT 27.160 30.670 27.520 31.035 ;
        RECT 27.600 30.670 27.960 31.035 ;
        RECT 28.040 30.670 28.400 31.035 ;
        RECT 28.480 30.670 28.840 31.035 ;
        RECT 55.160 30.670 55.520 31.035 ;
        RECT 55.600 30.670 55.960 31.035 ;
        RECT 56.040 30.670 56.400 31.035 ;
        RECT 56.480 30.670 56.840 31.035 ;
        RECT 83.160 30.670 83.520 31.035 ;
        RECT 83.600 30.670 83.960 31.035 ;
        RECT 84.040 30.670 84.400 31.035 ;
        RECT 84.480 30.670 84.840 31.035 ;
        RECT 111.160 24.020 111.520 24.385 ;
        RECT 111.600 24.020 111.960 24.385 ;
        RECT 112.040 24.020 112.400 24.385 ;
        RECT 112.480 24.020 112.840 24.385 ;
        RECT -0.840 22.620 -0.480 22.985 ;
        RECT -0.400 22.620 -0.040 22.985 ;
        RECT 0.040 22.620 0.400 22.985 ;
        RECT 0.480 22.620 0.840 22.985 ;
        RECT 27.160 -1.130 27.520 -0.765 ;
        RECT 27.600 -1.130 27.960 -0.765 ;
        RECT 28.040 -1.130 28.400 -0.765 ;
        RECT 28.480 -1.130 28.840 -0.765 ;
        RECT 55.160 -1.130 55.520 -0.765 ;
        RECT 55.600 -1.130 55.960 -0.765 ;
        RECT 56.040 -1.130 56.400 -0.765 ;
        RECT 56.480 -1.130 56.840 -0.765 ;
        RECT -0.800 -32.600 -0.400 -32.200 ;
        RECT -0.200 -32.600 0.200 -32.200 ;
        RECT 0.400 -32.600 0.800 -32.200 ;
        RECT 27.200 -32.600 27.600 -32.200 ;
        RECT 27.800 -32.600 28.200 -32.200 ;
        RECT 28.400 -32.600 28.800 -32.200 ;
        RECT 55.200 -32.600 55.600 -32.200 ;
        RECT 55.800 -32.600 56.200 -32.200 ;
        RECT 56.400 -32.600 56.800 -32.200 ;
        RECT 83.200 -32.600 83.600 -32.200 ;
        RECT 83.800 -32.600 84.200 -32.200 ;
        RECT 84.400 -32.600 84.800 -32.200 ;
        RECT 111.200 -32.600 111.600 -32.200 ;
        RECT 111.800 -32.600 112.200 -32.200 ;
        RECT 112.400 -32.600 112.800 -32.200 ;
        RECT -0.800 -33.200 -0.400 -32.800 ;
        RECT -0.200 -33.200 0.200 -32.800 ;
        RECT 0.400 -33.200 0.800 -32.800 ;
        RECT 27.200 -33.200 27.600 -32.800 ;
        RECT 27.800 -33.200 28.200 -32.800 ;
        RECT 28.400 -33.200 28.800 -32.800 ;
        RECT 55.200 -33.200 55.600 -32.800 ;
        RECT 55.800 -33.200 56.200 -32.800 ;
        RECT 56.400 -33.200 56.800 -32.800 ;
        RECT 83.200 -33.200 83.600 -32.800 ;
        RECT 83.800 -33.200 84.200 -32.800 ;
        RECT 84.400 -33.200 84.800 -32.800 ;
        RECT 111.200 -33.200 111.600 -32.800 ;
        RECT 111.800 -33.200 112.200 -32.800 ;
        RECT 112.400 -33.200 112.800 -32.800 ;
        RECT -0.800 -33.800 -0.400 -33.400 ;
        RECT -0.200 -33.800 0.200 -33.400 ;
        RECT 0.400 -33.800 0.800 -33.400 ;
        RECT 27.200 -33.800 27.600 -33.400 ;
        RECT 27.800 -33.800 28.200 -33.400 ;
        RECT 28.400 -33.800 28.800 -33.400 ;
        RECT 55.200 -33.800 55.600 -33.400 ;
        RECT 55.800 -33.800 56.200 -33.400 ;
        RECT 56.400 -33.800 56.800 -33.400 ;
        RECT 83.200 -33.800 83.600 -33.400 ;
        RECT 83.800 -33.800 84.200 -33.400 ;
        RECT 84.400 -33.800 84.800 -33.400 ;
        RECT 111.200 -33.800 111.600 -33.400 ;
        RECT 111.800 -33.800 112.200 -33.400 ;
        RECT 112.400 -33.800 112.800 -33.400 ;
      LAYER met4 ;
        RECT -1.000 -34.000 1.000 63.000 ;
        RECT 27.000 -34.000 29.000 63.000 ;
        RECT 55.000 -34.000 57.000 63.000 ;
        RECT 83.000 -34.000 85.000 63.000 ;
        RECT 111.000 -34.000 113.000 63.000 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 5.495 24.105 7.255 25.710 ;
      LAYER pwell ;
        RECT 2.180 23.585 3.985 23.815 ;
        RECT 1.695 22.905 3.985 23.585 ;
        RECT 1.840 22.715 2.010 22.905 ;
        RECT 5.830 22.715 6.000 22.885 ;
        RECT 10.980 15.470 100.050 22.570 ;
        RECT 103.000 20.000 106.000 25.000 ;
        RECT 103.000 19.000 111.000 20.000 ;
        RECT 105.000 17.000 111.000 19.000 ;
        RECT 2.500 7.270 109.280 14.370 ;
      LAYER li1 ;
        RECT 1.775 24.865 2.035 25.265 ;
        RECT 1.775 24.695 3.140 24.865 ;
        RECT 2.405 23.625 3.140 24.695 ;
        RECT 3.665 24.750 3.905 24.755 ;
        RECT 4.180 24.750 5.505 24.960 ;
        RECT 3.665 24.740 5.505 24.750 ;
        RECT 3.665 24.530 4.400 24.740 ;
        RECT 5.285 24.535 5.505 24.740 ;
        RECT 5.770 24.535 6.290 24.540 ;
        RECT 3.665 23.775 3.905 24.530 ;
        RECT 5.285 24.315 6.290 24.535 ;
        RECT 1.775 23.455 3.140 23.625 ;
        RECT 1.775 23.055 2.035 23.455 ;
        RECT 5.770 23.055 6.290 24.315 ;
        RECT 6.460 23.715 6.980 25.265 ;
        RECT 18.400 22.950 18.780 23.000 ;
        RECT 17.450 22.590 18.780 22.950 ;
        RECT 18.400 22.540 18.780 22.590 ;
        RECT 11.670 16.090 11.960 21.540 ;
        RECT 16.050 16.090 16.340 21.540 ;
        RECT 17.190 16.090 17.480 21.540 ;
        RECT 19.375 16.500 19.675 29.090 ;
        RECT 20.270 22.950 20.650 23.000 ;
        RECT 20.270 22.590 21.600 22.950 ;
        RECT 20.270 22.540 20.650 22.590 ;
        RECT 21.570 16.090 21.860 21.540 ;
        RECT 22.710 16.090 23.000 21.540 ;
        RECT 24.900 16.500 25.200 29.090 ;
        RECT 27.250 22.950 27.630 23.000 ;
        RECT 36.110 22.950 36.490 23.000 ;
        RECT 26.300 22.590 27.630 22.950 ;
        RECT 35.160 22.590 36.490 22.950 ;
        RECT 27.250 22.540 27.630 22.590 ;
        RECT 36.110 22.540 36.490 22.590 ;
        RECT 26.040 16.090 26.330 21.540 ;
        RECT 29.380 16.090 29.670 21.540 ;
        RECT 33.760 16.090 34.050 21.540 ;
        RECT 34.900 16.090 35.190 21.540 ;
        RECT 37.085 16.500 37.385 29.090 ;
        RECT 37.980 22.950 38.360 23.000 ;
        RECT 37.980 22.590 39.310 22.950 ;
        RECT 37.980 22.540 38.360 22.590 ;
        RECT 39.280 16.090 39.570 21.540 ;
        RECT 40.420 16.090 40.710 21.540 ;
        RECT 42.610 16.500 42.910 29.090 ;
        RECT 44.960 22.950 45.340 23.000 ;
        RECT 53.820 22.950 54.200 23.000 ;
        RECT 44.010 22.590 45.340 22.950 ;
        RECT 52.870 22.590 54.200 22.950 ;
        RECT 44.960 22.540 45.340 22.590 ;
        RECT 53.820 22.540 54.200 22.590 ;
        RECT 43.750 16.090 44.040 21.540 ;
        RECT 47.090 16.090 47.380 21.540 ;
        RECT 51.470 16.090 51.760 21.540 ;
        RECT 52.610 16.090 52.900 21.540 ;
        RECT 54.795 16.500 55.095 29.090 ;
        RECT 55.690 22.950 56.070 23.000 ;
        RECT 55.690 22.590 57.020 22.950 ;
        RECT 55.690 22.540 56.070 22.590 ;
        RECT 56.990 16.090 57.280 21.540 ;
        RECT 58.130 16.090 58.420 21.540 ;
        RECT 60.320 16.500 60.620 29.090 ;
        RECT 62.670 22.950 63.050 23.000 ;
        RECT 71.530 22.950 71.910 23.000 ;
        RECT 61.720 22.590 63.050 22.950 ;
        RECT 70.580 22.590 71.910 22.950 ;
        RECT 62.670 22.540 63.050 22.590 ;
        RECT 71.530 22.540 71.910 22.590 ;
        RECT 61.460 16.090 61.750 21.540 ;
        RECT 64.800 16.090 65.090 21.540 ;
        RECT 69.180 16.090 69.470 21.540 ;
        RECT 70.320 16.090 70.610 21.540 ;
        RECT 72.505 16.500 72.805 29.090 ;
        RECT 73.400 22.950 73.780 23.000 ;
        RECT 73.400 22.590 74.730 22.950 ;
        RECT 73.400 22.540 73.780 22.590 ;
        RECT 74.700 16.090 74.990 21.540 ;
        RECT 75.840 16.090 76.130 21.540 ;
        RECT 78.030 16.500 78.330 29.090 ;
        RECT 80.380 22.950 80.760 23.000 ;
        RECT 89.240 22.950 89.620 23.000 ;
        RECT 79.430 22.590 80.760 22.950 ;
        RECT 88.290 22.590 89.620 22.950 ;
        RECT 80.380 22.540 80.760 22.590 ;
        RECT 89.240 22.540 89.620 22.590 ;
        RECT 79.170 16.090 79.460 21.540 ;
        RECT 82.510 16.090 82.800 21.540 ;
        RECT 86.890 16.090 87.180 21.540 ;
        RECT 88.030 16.090 88.320 21.540 ;
        RECT 90.215 16.500 90.515 29.090 ;
        RECT 91.110 22.950 91.490 23.000 ;
        RECT 91.110 22.590 92.440 22.950 ;
        RECT 91.110 22.540 91.490 22.590 ;
        RECT 92.410 16.090 92.700 21.540 ;
        RECT 93.550 16.090 93.840 21.540 ;
        RECT 95.740 16.500 96.040 29.090 ;
        RECT 98.090 22.950 98.470 23.000 ;
        RECT 97.140 22.590 98.470 22.950 ;
        RECT 98.090 22.540 98.470 22.590 ;
        RECT 96.880 16.090 97.170 21.540 ;
        RECT 103.500 19.500 105.500 19.865 ;
        RECT 104.500 18.500 105.865 19.500 ;
        RECT 105.500 17.500 105.865 18.500 ;
        RECT 11.160 15.730 13.050 16.090 ;
        RECT 14.840 15.730 18.690 16.090 ;
        RECT 20.350 15.730 24.200 16.090 ;
        RECT 26.040 15.730 27.440 16.090 ;
        RECT 28.870 15.730 30.760 16.090 ;
        RECT 32.550 15.730 36.400 16.090 ;
        RECT 38.060 15.730 41.910 16.090 ;
        RECT 43.750 15.730 45.150 16.090 ;
        RECT 46.580 15.730 48.470 16.090 ;
        RECT 50.260 15.730 54.110 16.090 ;
        RECT 55.770 15.730 59.620 16.090 ;
        RECT 61.460 15.730 62.860 16.090 ;
        RECT 64.290 15.730 66.180 16.090 ;
        RECT 67.970 15.730 71.820 16.090 ;
        RECT 73.480 15.730 77.330 16.090 ;
        RECT 79.170 15.730 80.570 16.090 ;
        RECT 82.000 15.730 83.890 16.090 ;
        RECT 85.680 15.730 89.530 16.090 ;
        RECT 91.190 15.730 95.040 16.090 ;
        RECT 96.880 15.730 98.280 16.090 ;
        RECT 4.270 13.750 5.670 14.110 ;
        RECT 7.510 13.750 11.360 14.110 ;
        RECT 13.020 13.750 16.870 14.110 ;
        RECT 18.660 13.750 20.550 14.110 ;
        RECT 21.980 13.750 23.380 14.110 ;
        RECT 25.220 13.750 29.070 14.110 ;
        RECT 30.730 13.750 34.580 14.110 ;
        RECT 36.370 13.750 38.260 14.110 ;
        RECT 39.690 13.750 41.090 14.110 ;
        RECT 42.930 13.750 46.780 14.110 ;
        RECT 48.440 13.750 52.290 14.110 ;
        RECT 54.080 13.750 55.970 14.110 ;
        RECT 57.400 13.750 58.800 14.110 ;
        RECT 60.640 13.750 64.490 14.110 ;
        RECT 66.150 13.750 70.000 14.110 ;
        RECT 71.790 13.750 73.680 14.110 ;
        RECT 75.110 13.750 76.510 14.110 ;
        RECT 78.350 13.750 82.200 14.110 ;
        RECT 83.860 13.750 87.710 14.110 ;
        RECT 89.500 13.750 91.390 14.110 ;
        RECT 92.820 13.750 94.220 14.110 ;
        RECT 96.060 13.750 99.910 14.110 ;
        RECT 101.570 13.750 105.420 14.110 ;
        RECT 107.210 13.750 109.100 14.110 ;
        RECT 5.380 8.300 5.670 13.750 ;
        RECT 4.080 7.250 4.460 7.300 ;
        RECT 4.080 6.890 5.410 7.250 ;
        RECT 4.080 6.840 4.460 6.890 ;
        RECT 6.510 0.750 6.810 13.340 ;
        RECT 8.710 8.300 9.000 13.750 ;
        RECT 9.850 8.300 10.140 13.750 ;
        RECT 11.060 7.250 11.440 7.300 ;
        RECT 10.110 6.890 11.440 7.250 ;
        RECT 11.060 6.840 11.440 6.890 ;
        RECT 12.035 0.750 12.335 13.340 ;
        RECT 14.230 8.300 14.520 13.750 ;
        RECT 15.370 8.300 15.660 13.750 ;
        RECT 19.750 8.300 20.040 13.750 ;
        RECT 23.090 8.300 23.380 13.750 ;
        RECT 12.930 7.250 13.310 7.300 ;
        RECT 21.790 7.250 22.170 7.300 ;
        RECT 12.930 6.890 14.260 7.250 ;
        RECT 21.790 6.890 23.120 7.250 ;
        RECT 12.930 6.840 13.310 6.890 ;
        RECT 21.790 6.840 22.170 6.890 ;
        RECT 24.220 0.750 24.520 13.340 ;
        RECT 26.420 8.300 26.710 13.750 ;
        RECT 27.560 8.300 27.850 13.750 ;
        RECT 28.770 7.250 29.150 7.300 ;
        RECT 27.820 6.890 29.150 7.250 ;
        RECT 28.770 6.840 29.150 6.890 ;
        RECT 29.745 0.750 30.045 13.340 ;
        RECT 31.940 8.300 32.230 13.750 ;
        RECT 33.080 8.300 33.370 13.750 ;
        RECT 37.460 8.300 37.750 13.750 ;
        RECT 40.800 8.300 41.090 13.750 ;
        RECT 30.640 7.250 31.020 7.300 ;
        RECT 39.500 7.250 39.880 7.300 ;
        RECT 30.640 6.890 31.970 7.250 ;
        RECT 39.500 6.890 40.830 7.250 ;
        RECT 30.640 6.840 31.020 6.890 ;
        RECT 39.500 6.840 39.880 6.890 ;
        RECT 41.930 0.750 42.230 13.340 ;
        RECT 44.130 8.300 44.420 13.750 ;
        RECT 45.270 8.300 45.560 13.750 ;
        RECT 46.480 7.250 46.860 7.300 ;
        RECT 45.530 6.890 46.860 7.250 ;
        RECT 46.480 6.840 46.860 6.890 ;
        RECT 47.455 0.750 47.755 13.340 ;
        RECT 49.650 8.300 49.940 13.750 ;
        RECT 50.790 8.300 51.080 13.750 ;
        RECT 55.170 8.300 55.460 13.750 ;
        RECT 58.510 8.300 58.800 13.750 ;
        RECT 48.350 7.250 48.730 7.300 ;
        RECT 57.210 7.250 57.590 7.300 ;
        RECT 48.350 6.890 49.680 7.250 ;
        RECT 57.210 6.890 58.540 7.250 ;
        RECT 48.350 6.840 48.730 6.890 ;
        RECT 57.210 6.840 57.590 6.890 ;
        RECT 59.640 0.750 59.940 13.340 ;
        RECT 61.840 8.300 62.130 13.750 ;
        RECT 62.980 8.300 63.270 13.750 ;
        RECT 64.190 7.250 64.570 7.300 ;
        RECT 63.240 6.890 64.570 7.250 ;
        RECT 64.190 6.840 64.570 6.890 ;
        RECT 65.165 0.750 65.465 13.340 ;
        RECT 67.360 8.300 67.650 13.750 ;
        RECT 68.500 8.300 68.790 13.750 ;
        RECT 72.880 8.300 73.170 13.750 ;
        RECT 76.220 8.300 76.510 13.750 ;
        RECT 66.060 7.250 66.440 7.300 ;
        RECT 74.920 7.250 75.300 7.300 ;
        RECT 66.060 6.890 67.390 7.250 ;
        RECT 74.920 6.890 76.250 7.250 ;
        RECT 66.060 6.840 66.440 6.890 ;
        RECT 74.920 6.840 75.300 6.890 ;
        RECT 77.350 0.750 77.650 13.340 ;
        RECT 79.550 8.300 79.840 13.750 ;
        RECT 80.690 8.300 80.980 13.750 ;
        RECT 81.900 7.250 82.280 7.300 ;
        RECT 80.950 6.890 82.280 7.250 ;
        RECT 81.900 6.840 82.280 6.890 ;
        RECT 82.875 0.750 83.175 13.340 ;
        RECT 85.070 8.300 85.360 13.750 ;
        RECT 86.210 8.300 86.500 13.750 ;
        RECT 90.590 8.300 90.880 13.750 ;
        RECT 93.930 8.300 94.220 13.750 ;
        RECT 83.770 7.250 84.150 7.300 ;
        RECT 92.630 7.250 93.010 7.300 ;
        RECT 83.770 6.890 85.100 7.250 ;
        RECT 92.630 6.890 93.960 7.250 ;
        RECT 83.770 6.840 84.150 6.890 ;
        RECT 92.630 6.840 93.010 6.890 ;
        RECT 95.060 0.750 95.360 13.340 ;
        RECT 97.260 8.300 97.550 13.750 ;
        RECT 98.400 8.300 98.690 13.750 ;
        RECT 99.610 7.250 99.990 7.300 ;
        RECT 98.660 6.890 99.990 7.250 ;
        RECT 99.610 6.840 99.990 6.890 ;
        RECT 100.585 0.750 100.885 13.340 ;
        RECT 102.780 8.300 103.070 13.750 ;
        RECT 103.920 8.300 104.210 13.750 ;
        RECT 108.300 8.300 108.590 13.750 ;
        RECT 101.480 7.250 101.860 7.300 ;
        RECT 101.480 6.890 102.810 7.250 ;
        RECT 101.480 6.840 101.860 6.890 ;
      LAYER mcon ;
        RECT 17.450 22.620 17.750 22.920 ;
        RECT 17.940 22.620 18.240 22.920 ;
        RECT 18.430 22.620 18.730 22.920 ;
        RECT 20.320 22.620 20.620 22.920 ;
        RECT 20.810 22.620 21.110 22.920 ;
        RECT 21.300 22.620 21.600 22.920 ;
        RECT 19.375 21.260 19.675 21.560 ;
        RECT 26.300 22.620 26.600 22.920 ;
        RECT 26.790 22.620 27.090 22.920 ;
        RECT 27.280 22.620 27.580 22.920 ;
        RECT 35.160 22.620 35.460 22.920 ;
        RECT 35.650 22.620 35.950 22.920 ;
        RECT 36.140 22.620 36.440 22.920 ;
        RECT 24.900 21.260 25.200 21.560 ;
        RECT 38.030 22.620 38.330 22.920 ;
        RECT 38.520 22.620 38.820 22.920 ;
        RECT 39.010 22.620 39.310 22.920 ;
        RECT 37.085 21.260 37.385 21.560 ;
        RECT 44.010 22.620 44.310 22.920 ;
        RECT 44.500 22.620 44.800 22.920 ;
        RECT 44.990 22.620 45.290 22.920 ;
        RECT 52.870 22.620 53.170 22.920 ;
        RECT 53.360 22.620 53.660 22.920 ;
        RECT 53.850 22.620 54.150 22.920 ;
        RECT 42.610 21.260 42.910 21.560 ;
        RECT 55.740 22.620 56.040 22.920 ;
        RECT 56.230 22.620 56.530 22.920 ;
        RECT 56.720 22.620 57.020 22.920 ;
        RECT 54.795 21.260 55.095 21.560 ;
        RECT 61.720 22.620 62.020 22.920 ;
        RECT 62.210 22.620 62.510 22.920 ;
        RECT 62.700 22.620 63.000 22.920 ;
        RECT 70.580 22.620 70.880 22.920 ;
        RECT 71.070 22.620 71.370 22.920 ;
        RECT 71.560 22.620 71.860 22.920 ;
        RECT 60.320 21.260 60.620 21.560 ;
        RECT 73.450 22.620 73.750 22.920 ;
        RECT 73.940 22.620 74.240 22.920 ;
        RECT 74.430 22.620 74.730 22.920 ;
        RECT 72.505 21.260 72.805 21.560 ;
        RECT 79.430 22.620 79.730 22.920 ;
        RECT 79.920 22.620 80.220 22.920 ;
        RECT 80.410 22.620 80.710 22.920 ;
        RECT 88.290 22.620 88.590 22.920 ;
        RECT 88.780 22.620 89.080 22.920 ;
        RECT 89.270 22.620 89.570 22.920 ;
        RECT 78.030 21.260 78.330 21.560 ;
        RECT 91.160 22.620 91.460 22.920 ;
        RECT 91.650 22.620 91.950 22.920 ;
        RECT 92.140 22.620 92.440 22.920 ;
        RECT 90.215 21.260 90.515 21.560 ;
        RECT 97.140 22.620 97.440 22.920 ;
        RECT 97.630 22.620 97.930 22.920 ;
        RECT 98.120 22.620 98.420 22.920 ;
        RECT 95.740 21.260 96.040 21.560 ;
        RECT 104.590 19.120 104.890 19.420 ;
        RECT 105.110 19.120 105.410 19.420 ;
        RECT 104.590 18.600 104.890 18.900 ;
        RECT 105.110 18.600 105.410 18.900 ;
        RECT 11.220 15.760 11.520 16.060 ;
        RECT 11.710 15.760 12.010 16.060 ;
        RECT 12.200 15.760 12.500 16.060 ;
        RECT 12.690 15.760 12.990 16.060 ;
        RECT 14.900 15.760 15.200 16.060 ;
        RECT 15.390 15.760 15.690 16.060 ;
        RECT 15.880 15.760 16.180 16.060 ;
        RECT 16.370 15.760 16.670 16.060 ;
        RECT 16.860 15.760 17.160 16.060 ;
        RECT 17.350 15.760 17.650 16.060 ;
        RECT 17.840 15.760 18.140 16.060 ;
        RECT 18.330 15.760 18.630 16.060 ;
        RECT 20.410 15.760 20.710 16.060 ;
        RECT 20.900 15.760 21.200 16.060 ;
        RECT 21.390 15.760 21.690 16.060 ;
        RECT 21.880 15.760 22.180 16.060 ;
        RECT 22.370 15.760 22.670 16.060 ;
        RECT 22.860 15.760 23.160 16.060 ;
        RECT 23.350 15.760 23.650 16.060 ;
        RECT 23.840 15.760 24.140 16.060 ;
        RECT 26.100 15.760 26.400 16.060 ;
        RECT 26.590 15.760 26.890 16.060 ;
        RECT 27.080 15.760 27.380 16.060 ;
        RECT 28.930 15.760 29.230 16.060 ;
        RECT 29.420 15.760 29.720 16.060 ;
        RECT 29.910 15.760 30.210 16.060 ;
        RECT 30.400 15.760 30.700 16.060 ;
        RECT 32.610 15.760 32.910 16.060 ;
        RECT 33.100 15.760 33.400 16.060 ;
        RECT 33.590 15.760 33.890 16.060 ;
        RECT 34.080 15.760 34.380 16.060 ;
        RECT 34.570 15.760 34.870 16.060 ;
        RECT 35.060 15.760 35.360 16.060 ;
        RECT 35.550 15.760 35.850 16.060 ;
        RECT 36.040 15.760 36.340 16.060 ;
        RECT 38.120 15.760 38.420 16.060 ;
        RECT 38.610 15.760 38.910 16.060 ;
        RECT 39.100 15.760 39.400 16.060 ;
        RECT 39.590 15.760 39.890 16.060 ;
        RECT 40.080 15.760 40.380 16.060 ;
        RECT 40.570 15.760 40.870 16.060 ;
        RECT 41.060 15.760 41.360 16.060 ;
        RECT 41.550 15.760 41.850 16.060 ;
        RECT 43.810 15.760 44.110 16.060 ;
        RECT 44.300 15.760 44.600 16.060 ;
        RECT 44.790 15.760 45.090 16.060 ;
        RECT 46.640 15.760 46.940 16.060 ;
        RECT 47.130 15.760 47.430 16.060 ;
        RECT 47.620 15.760 47.920 16.060 ;
        RECT 48.110 15.760 48.410 16.060 ;
        RECT 50.320 15.760 50.620 16.060 ;
        RECT 50.810 15.760 51.110 16.060 ;
        RECT 51.300 15.760 51.600 16.060 ;
        RECT 51.790 15.760 52.090 16.060 ;
        RECT 52.280 15.760 52.580 16.060 ;
        RECT 52.770 15.760 53.070 16.060 ;
        RECT 53.260 15.760 53.560 16.060 ;
        RECT 53.750 15.760 54.050 16.060 ;
        RECT 55.830 15.760 56.130 16.060 ;
        RECT 56.320 15.760 56.620 16.060 ;
        RECT 56.810 15.760 57.110 16.060 ;
        RECT 57.300 15.760 57.600 16.060 ;
        RECT 57.790 15.760 58.090 16.060 ;
        RECT 58.280 15.760 58.580 16.060 ;
        RECT 58.770 15.760 59.070 16.060 ;
        RECT 59.260 15.760 59.560 16.060 ;
        RECT 61.520 15.760 61.820 16.060 ;
        RECT 62.010 15.760 62.310 16.060 ;
        RECT 62.500 15.760 62.800 16.060 ;
        RECT 64.350 15.760 64.650 16.060 ;
        RECT 64.840 15.760 65.140 16.060 ;
        RECT 65.330 15.760 65.630 16.060 ;
        RECT 65.820 15.760 66.120 16.060 ;
        RECT 68.030 15.760 68.330 16.060 ;
        RECT 68.520 15.760 68.820 16.060 ;
        RECT 69.010 15.760 69.310 16.060 ;
        RECT 69.500 15.760 69.800 16.060 ;
        RECT 69.990 15.760 70.290 16.060 ;
        RECT 70.480 15.760 70.780 16.060 ;
        RECT 70.970 15.760 71.270 16.060 ;
        RECT 71.460 15.760 71.760 16.060 ;
        RECT 73.540 15.760 73.840 16.060 ;
        RECT 74.030 15.760 74.330 16.060 ;
        RECT 74.520 15.760 74.820 16.060 ;
        RECT 75.010 15.760 75.310 16.060 ;
        RECT 75.500 15.760 75.800 16.060 ;
        RECT 75.990 15.760 76.290 16.060 ;
        RECT 76.480 15.760 76.780 16.060 ;
        RECT 76.970 15.760 77.270 16.060 ;
        RECT 79.230 15.760 79.530 16.060 ;
        RECT 79.720 15.760 80.020 16.060 ;
        RECT 80.210 15.760 80.510 16.060 ;
        RECT 82.060 15.760 82.360 16.060 ;
        RECT 82.550 15.760 82.850 16.060 ;
        RECT 83.040 15.760 83.340 16.060 ;
        RECT 83.530 15.760 83.830 16.060 ;
        RECT 85.740 15.760 86.040 16.060 ;
        RECT 86.230 15.760 86.530 16.060 ;
        RECT 86.720 15.760 87.020 16.060 ;
        RECT 87.210 15.760 87.510 16.060 ;
        RECT 87.700 15.760 88.000 16.060 ;
        RECT 88.190 15.760 88.490 16.060 ;
        RECT 88.680 15.760 88.980 16.060 ;
        RECT 89.170 15.760 89.470 16.060 ;
        RECT 91.250 15.760 91.550 16.060 ;
        RECT 91.740 15.760 92.040 16.060 ;
        RECT 92.230 15.760 92.530 16.060 ;
        RECT 92.720 15.760 93.020 16.060 ;
        RECT 93.210 15.760 93.510 16.060 ;
        RECT 93.700 15.760 94.000 16.060 ;
        RECT 94.190 15.760 94.490 16.060 ;
        RECT 94.680 15.760 94.980 16.060 ;
        RECT 96.940 15.760 97.240 16.060 ;
        RECT 97.430 15.760 97.730 16.060 ;
        RECT 97.920 15.760 98.220 16.060 ;
        RECT 4.330 13.780 4.630 14.080 ;
        RECT 4.820 13.780 5.120 14.080 ;
        RECT 5.310 13.780 5.610 14.080 ;
        RECT 7.570 13.780 7.870 14.080 ;
        RECT 8.060 13.780 8.360 14.080 ;
        RECT 8.550 13.780 8.850 14.080 ;
        RECT 9.040 13.780 9.340 14.080 ;
        RECT 9.530 13.780 9.830 14.080 ;
        RECT 10.020 13.780 10.320 14.080 ;
        RECT 10.510 13.780 10.810 14.080 ;
        RECT 11.000 13.780 11.300 14.080 ;
        RECT 13.080 13.780 13.380 14.080 ;
        RECT 13.570 13.780 13.870 14.080 ;
        RECT 14.060 13.780 14.360 14.080 ;
        RECT 14.550 13.780 14.850 14.080 ;
        RECT 15.040 13.780 15.340 14.080 ;
        RECT 15.530 13.780 15.830 14.080 ;
        RECT 16.020 13.780 16.320 14.080 ;
        RECT 16.510 13.780 16.810 14.080 ;
        RECT 18.720 13.780 19.020 14.080 ;
        RECT 19.210 13.780 19.510 14.080 ;
        RECT 19.700 13.780 20.000 14.080 ;
        RECT 20.190 13.780 20.490 14.080 ;
        RECT 22.040 13.780 22.340 14.080 ;
        RECT 22.530 13.780 22.830 14.080 ;
        RECT 23.020 13.780 23.320 14.080 ;
        RECT 25.280 13.780 25.580 14.080 ;
        RECT 25.770 13.780 26.070 14.080 ;
        RECT 26.260 13.780 26.560 14.080 ;
        RECT 26.750 13.780 27.050 14.080 ;
        RECT 27.240 13.780 27.540 14.080 ;
        RECT 27.730 13.780 28.030 14.080 ;
        RECT 28.220 13.780 28.520 14.080 ;
        RECT 28.710 13.780 29.010 14.080 ;
        RECT 30.790 13.780 31.090 14.080 ;
        RECT 31.280 13.780 31.580 14.080 ;
        RECT 31.770 13.780 32.070 14.080 ;
        RECT 32.260 13.780 32.560 14.080 ;
        RECT 32.750 13.780 33.050 14.080 ;
        RECT 33.240 13.780 33.540 14.080 ;
        RECT 33.730 13.780 34.030 14.080 ;
        RECT 34.220 13.780 34.520 14.080 ;
        RECT 36.430 13.780 36.730 14.080 ;
        RECT 36.920 13.780 37.220 14.080 ;
        RECT 37.410 13.780 37.710 14.080 ;
        RECT 37.900 13.780 38.200 14.080 ;
        RECT 39.750 13.780 40.050 14.080 ;
        RECT 40.240 13.780 40.540 14.080 ;
        RECT 40.730 13.780 41.030 14.080 ;
        RECT 42.990 13.780 43.290 14.080 ;
        RECT 43.480 13.780 43.780 14.080 ;
        RECT 43.970 13.780 44.270 14.080 ;
        RECT 44.460 13.780 44.760 14.080 ;
        RECT 44.950 13.780 45.250 14.080 ;
        RECT 45.440 13.780 45.740 14.080 ;
        RECT 45.930 13.780 46.230 14.080 ;
        RECT 46.420 13.780 46.720 14.080 ;
        RECT 48.500 13.780 48.800 14.080 ;
        RECT 48.990 13.780 49.290 14.080 ;
        RECT 49.480 13.780 49.780 14.080 ;
        RECT 49.970 13.780 50.270 14.080 ;
        RECT 50.460 13.780 50.760 14.080 ;
        RECT 50.950 13.780 51.250 14.080 ;
        RECT 51.440 13.780 51.740 14.080 ;
        RECT 51.930 13.780 52.230 14.080 ;
        RECT 54.140 13.780 54.440 14.080 ;
        RECT 54.630 13.780 54.930 14.080 ;
        RECT 55.120 13.780 55.420 14.080 ;
        RECT 55.610 13.780 55.910 14.080 ;
        RECT 57.460 13.780 57.760 14.080 ;
        RECT 57.950 13.780 58.250 14.080 ;
        RECT 58.440 13.780 58.740 14.080 ;
        RECT 60.700 13.780 61.000 14.080 ;
        RECT 61.190 13.780 61.490 14.080 ;
        RECT 61.680 13.780 61.980 14.080 ;
        RECT 62.170 13.780 62.470 14.080 ;
        RECT 62.660 13.780 62.960 14.080 ;
        RECT 63.150 13.780 63.450 14.080 ;
        RECT 63.640 13.780 63.940 14.080 ;
        RECT 64.130 13.780 64.430 14.080 ;
        RECT 66.210 13.780 66.510 14.080 ;
        RECT 66.700 13.780 67.000 14.080 ;
        RECT 67.190 13.780 67.490 14.080 ;
        RECT 67.680 13.780 67.980 14.080 ;
        RECT 68.170 13.780 68.470 14.080 ;
        RECT 68.660 13.780 68.960 14.080 ;
        RECT 69.150 13.780 69.450 14.080 ;
        RECT 69.640 13.780 69.940 14.080 ;
        RECT 71.850 13.780 72.150 14.080 ;
        RECT 72.340 13.780 72.640 14.080 ;
        RECT 72.830 13.780 73.130 14.080 ;
        RECT 73.320 13.780 73.620 14.080 ;
        RECT 75.170 13.780 75.470 14.080 ;
        RECT 75.660 13.780 75.960 14.080 ;
        RECT 76.150 13.780 76.450 14.080 ;
        RECT 78.410 13.780 78.710 14.080 ;
        RECT 78.900 13.780 79.200 14.080 ;
        RECT 79.390 13.780 79.690 14.080 ;
        RECT 79.880 13.780 80.180 14.080 ;
        RECT 80.370 13.780 80.670 14.080 ;
        RECT 80.860 13.780 81.160 14.080 ;
        RECT 81.350 13.780 81.650 14.080 ;
        RECT 81.840 13.780 82.140 14.080 ;
        RECT 83.920 13.780 84.220 14.080 ;
        RECT 84.410 13.780 84.710 14.080 ;
        RECT 84.900 13.780 85.200 14.080 ;
        RECT 85.390 13.780 85.690 14.080 ;
        RECT 85.880 13.780 86.180 14.080 ;
        RECT 86.370 13.780 86.670 14.080 ;
        RECT 86.860 13.780 87.160 14.080 ;
        RECT 87.350 13.780 87.650 14.080 ;
        RECT 89.560 13.780 89.860 14.080 ;
        RECT 90.050 13.780 90.350 14.080 ;
        RECT 90.540 13.780 90.840 14.080 ;
        RECT 91.030 13.780 91.330 14.080 ;
        RECT 92.880 13.780 93.180 14.080 ;
        RECT 93.370 13.780 93.670 14.080 ;
        RECT 93.860 13.780 94.160 14.080 ;
        RECT 96.120 13.780 96.420 14.080 ;
        RECT 96.610 13.780 96.910 14.080 ;
        RECT 97.100 13.780 97.400 14.080 ;
        RECT 97.590 13.780 97.890 14.080 ;
        RECT 98.080 13.780 98.380 14.080 ;
        RECT 98.570 13.780 98.870 14.080 ;
        RECT 99.060 13.780 99.360 14.080 ;
        RECT 99.550 13.780 99.850 14.080 ;
        RECT 101.630 13.780 101.930 14.080 ;
        RECT 102.120 13.780 102.420 14.080 ;
        RECT 102.610 13.780 102.910 14.080 ;
        RECT 103.100 13.780 103.400 14.080 ;
        RECT 103.590 13.780 103.890 14.080 ;
        RECT 104.080 13.780 104.380 14.080 ;
        RECT 104.570 13.780 104.870 14.080 ;
        RECT 105.060 13.780 105.360 14.080 ;
        RECT 107.270 13.780 107.570 14.080 ;
        RECT 107.760 13.780 108.060 14.080 ;
        RECT 108.250 13.780 108.550 14.080 ;
        RECT 108.740 13.780 109.040 14.080 ;
        RECT 6.510 8.280 6.810 8.580 ;
        RECT 4.130 6.920 4.430 7.220 ;
        RECT 4.620 6.920 4.920 7.220 ;
        RECT 5.110 6.920 5.410 7.220 ;
        RECT 12.035 8.280 12.335 8.580 ;
        RECT 10.110 6.920 10.410 7.220 ;
        RECT 10.600 6.920 10.900 7.220 ;
        RECT 11.090 6.920 11.390 7.220 ;
        RECT 24.220 8.280 24.520 8.580 ;
        RECT 12.980 6.920 13.280 7.220 ;
        RECT 13.470 6.920 13.770 7.220 ;
        RECT 13.960 6.920 14.260 7.220 ;
        RECT 21.840 6.920 22.140 7.220 ;
        RECT 22.330 6.920 22.630 7.220 ;
        RECT 22.820 6.920 23.120 7.220 ;
        RECT 29.745 8.280 30.045 8.580 ;
        RECT 27.820 6.920 28.120 7.220 ;
        RECT 28.310 6.920 28.610 7.220 ;
        RECT 28.800 6.920 29.100 7.220 ;
        RECT 41.930 8.280 42.230 8.580 ;
        RECT 30.690 6.920 30.990 7.220 ;
        RECT 31.180 6.920 31.480 7.220 ;
        RECT 31.670 6.920 31.970 7.220 ;
        RECT 39.550 6.920 39.850 7.220 ;
        RECT 40.040 6.920 40.340 7.220 ;
        RECT 40.530 6.920 40.830 7.220 ;
        RECT 47.455 8.280 47.755 8.580 ;
        RECT 45.530 6.920 45.830 7.220 ;
        RECT 46.020 6.920 46.320 7.220 ;
        RECT 46.510 6.920 46.810 7.220 ;
        RECT 59.640 8.280 59.940 8.580 ;
        RECT 48.400 6.920 48.700 7.220 ;
        RECT 48.890 6.920 49.190 7.220 ;
        RECT 49.380 6.920 49.680 7.220 ;
        RECT 57.260 6.920 57.560 7.220 ;
        RECT 57.750 6.920 58.050 7.220 ;
        RECT 58.240 6.920 58.540 7.220 ;
        RECT 65.165 8.280 65.465 8.580 ;
        RECT 63.240 6.920 63.540 7.220 ;
        RECT 63.730 6.920 64.030 7.220 ;
        RECT 64.220 6.920 64.520 7.220 ;
        RECT 77.350 8.280 77.650 8.580 ;
        RECT 66.110 6.920 66.410 7.220 ;
        RECT 66.600 6.920 66.900 7.220 ;
        RECT 67.090 6.920 67.390 7.220 ;
        RECT 74.970 6.920 75.270 7.220 ;
        RECT 75.460 6.920 75.760 7.220 ;
        RECT 75.950 6.920 76.250 7.220 ;
        RECT 82.875 8.280 83.175 8.580 ;
        RECT 80.950 6.920 81.250 7.220 ;
        RECT 81.440 6.920 81.740 7.220 ;
        RECT 81.930 6.920 82.230 7.220 ;
        RECT 95.060 8.280 95.360 8.580 ;
        RECT 83.820 6.920 84.120 7.220 ;
        RECT 84.310 6.920 84.610 7.220 ;
        RECT 84.800 6.920 85.100 7.220 ;
        RECT 92.680 6.920 92.980 7.220 ;
        RECT 93.170 6.920 93.470 7.220 ;
        RECT 93.660 6.920 93.960 7.220 ;
        RECT 100.585 8.280 100.885 8.580 ;
        RECT 98.660 6.920 98.960 7.220 ;
        RECT 99.150 6.920 99.450 7.220 ;
        RECT 99.640 6.920 99.940 7.220 ;
        RECT 101.530 6.920 101.830 7.220 ;
        RECT 102.020 6.920 102.320 7.220 ;
        RECT 102.510 6.920 102.810 7.220 ;
      LAYER met1 ;
        RECT 17.390 22.590 21.660 22.950 ;
        RECT 26.240 22.590 27.740 22.950 ;
        RECT 35.100 22.590 39.370 22.950 ;
        RECT 43.950 22.590 45.450 22.950 ;
        RECT 52.810 22.590 57.080 22.950 ;
        RECT 61.660 22.590 63.160 22.950 ;
        RECT 70.520 22.590 74.790 22.950 ;
        RECT 79.370 22.590 80.870 22.950 ;
        RECT 88.230 22.590 92.500 22.950 ;
        RECT 97.080 22.590 98.580 22.950 ;
        RECT 18.005 21.590 18.365 22.590 ;
        RECT 26.790 21.590 27.150 22.590 ;
        RECT 35.715 21.590 36.075 22.590 ;
        RECT 44.500 21.590 44.860 22.590 ;
        RECT 53.425 21.590 53.785 22.590 ;
        RECT 62.210 21.590 62.570 22.590 ;
        RECT 71.135 21.590 71.495 22.590 ;
        RECT 79.920 21.590 80.280 22.590 ;
        RECT 88.845 21.590 89.205 22.590 ;
        RECT 97.630 21.590 97.990 22.590 ;
        RECT 9.620 21.230 18.365 21.590 ;
        RECT 19.315 21.230 36.075 21.590 ;
        RECT 37.025 21.230 53.785 21.590 ;
        RECT 54.735 21.230 71.495 21.590 ;
        RECT 72.445 21.230 89.205 21.590 ;
        RECT 90.155 21.230 101.360 21.590 ;
        RECT 9.620 16.000 9.980 21.230 ;
        RECT 1.350 15.640 9.980 16.000 ;
        RECT 10.980 15.670 100.050 16.150 ;
        RECT 101.000 16.000 101.360 21.230 ;
        RECT 104.500 18.500 105.500 19.515 ;
        RECT 101.000 15.640 110.500 16.000 ;
        RECT 1.350 8.610 1.710 15.640 ;
        RECT 2.500 13.690 109.280 14.170 ;
        RECT 110.140 8.610 110.500 15.640 ;
        RECT 1.350 8.250 12.395 8.610 ;
        RECT 13.345 8.250 30.105 8.610 ;
        RECT 31.055 8.250 47.815 8.610 ;
        RECT 48.765 8.250 65.525 8.610 ;
        RECT 66.475 8.250 83.235 8.610 ;
        RECT 84.185 8.250 100.945 8.610 ;
        RECT 101.895 8.250 110.500 8.610 ;
        RECT 4.560 7.250 4.920 8.250 ;
        RECT 13.345 7.250 13.705 8.250 ;
        RECT 22.270 7.250 22.630 8.250 ;
        RECT 31.055 7.250 31.415 8.250 ;
        RECT 39.980 7.250 40.340 8.250 ;
        RECT 48.765 7.250 49.125 8.250 ;
        RECT 57.690 7.250 58.050 8.250 ;
        RECT 66.475 7.250 66.835 8.250 ;
        RECT 75.400 7.250 75.760 8.250 ;
        RECT 84.185 7.250 84.545 8.250 ;
        RECT 93.110 7.250 93.470 8.250 ;
        RECT 101.895 7.250 102.255 8.250 ;
        RECT 3.970 6.890 5.470 7.250 ;
        RECT 10.050 6.890 14.320 7.250 ;
        RECT 21.680 6.890 23.180 7.250 ;
        RECT 27.760 6.890 32.030 7.250 ;
        RECT 39.390 6.890 40.890 7.250 ;
        RECT 45.470 6.890 49.740 7.250 ;
        RECT 57.100 6.890 58.600 7.250 ;
        RECT 63.180 6.890 67.450 7.250 ;
        RECT 74.810 6.890 76.310 7.250 ;
        RECT 80.890 6.890 85.160 7.250 ;
        RECT 92.520 6.890 94.020 7.250 ;
        RECT 98.600 6.890 102.870 7.250 ;
      LAYER via ;
        RECT 14.500 15.770 14.760 16.030 ;
        RECT 14.870 15.770 15.130 16.030 ;
        RECT 15.240 15.770 15.500 16.030 ;
        RECT 20.500 15.770 20.760 16.030 ;
        RECT 20.870 15.770 21.130 16.030 ;
        RECT 21.240 15.770 21.500 16.030 ;
        RECT 26.500 15.770 26.760 16.030 ;
        RECT 26.870 15.770 27.130 16.030 ;
        RECT 27.240 15.770 27.500 16.030 ;
        RECT 32.500 15.770 32.760 16.030 ;
        RECT 32.870 15.770 33.130 16.030 ;
        RECT 33.240 15.770 33.500 16.030 ;
        RECT 38.500 15.770 38.760 16.030 ;
        RECT 38.870 15.770 39.130 16.030 ;
        RECT 39.240 15.770 39.500 16.030 ;
        RECT 44.500 15.770 44.760 16.030 ;
        RECT 44.870 15.770 45.130 16.030 ;
        RECT 45.240 15.770 45.500 16.030 ;
        RECT 50.500 15.770 50.760 16.030 ;
        RECT 50.870 15.770 51.130 16.030 ;
        RECT 51.240 15.770 51.500 16.030 ;
        RECT 56.500 15.770 56.760 16.030 ;
        RECT 56.870 15.770 57.130 16.030 ;
        RECT 57.240 15.770 57.500 16.030 ;
        RECT 62.500 15.770 62.760 16.030 ;
        RECT 62.870 15.770 63.130 16.030 ;
        RECT 63.240 15.770 63.500 16.030 ;
        RECT 68.500 15.770 68.760 16.030 ;
        RECT 68.870 15.770 69.130 16.030 ;
        RECT 69.240 15.770 69.500 16.030 ;
        RECT 74.500 15.770 74.760 16.030 ;
        RECT 74.870 15.770 75.130 16.030 ;
        RECT 75.240 15.770 75.500 16.030 ;
        RECT 80.500 15.770 80.760 16.030 ;
        RECT 80.870 15.770 81.130 16.030 ;
        RECT 81.240 15.770 81.500 16.030 ;
        RECT 86.500 15.770 86.760 16.030 ;
        RECT 86.870 15.770 87.130 16.030 ;
        RECT 87.240 15.770 87.500 16.030 ;
        RECT 92.500 15.770 92.760 16.030 ;
        RECT 92.870 15.770 93.130 16.030 ;
        RECT 93.240 15.770 93.500 16.030 ;
        RECT 98.500 15.770 98.760 16.030 ;
        RECT 98.870 15.770 99.130 16.030 ;
        RECT 99.240 15.770 99.500 16.030 ;
        RECT 104.570 19.100 104.910 19.440 ;
        RECT 105.090 19.100 105.430 19.440 ;
        RECT 104.570 18.580 104.910 18.920 ;
        RECT 105.090 18.580 105.430 18.920 ;
        RECT 2.500 13.790 2.760 14.050 ;
        RECT 2.870 13.790 3.130 14.050 ;
        RECT 3.240 13.790 3.500 14.050 ;
        RECT 8.500 13.790 8.760 14.050 ;
        RECT 8.870 13.790 9.130 14.050 ;
        RECT 9.240 13.790 9.500 14.050 ;
        RECT 14.500 13.790 14.760 14.050 ;
        RECT 14.870 13.790 15.130 14.050 ;
        RECT 15.240 13.790 15.500 14.050 ;
        RECT 20.500 13.790 20.760 14.050 ;
        RECT 20.870 13.790 21.130 14.050 ;
        RECT 21.240 13.790 21.500 14.050 ;
        RECT 26.500 13.790 26.760 14.050 ;
        RECT 26.870 13.790 27.130 14.050 ;
        RECT 27.240 13.790 27.500 14.050 ;
        RECT 32.500 13.790 32.760 14.050 ;
        RECT 32.870 13.790 33.130 14.050 ;
        RECT 33.240 13.790 33.500 14.050 ;
        RECT 38.500 13.790 38.760 14.050 ;
        RECT 38.870 13.790 39.130 14.050 ;
        RECT 39.240 13.790 39.500 14.050 ;
        RECT 44.500 13.790 44.760 14.050 ;
        RECT 44.870 13.790 45.130 14.050 ;
        RECT 45.240 13.790 45.500 14.050 ;
        RECT 50.500 13.790 50.760 14.050 ;
        RECT 50.870 13.790 51.130 14.050 ;
        RECT 51.240 13.790 51.500 14.050 ;
        RECT 56.500 13.790 56.760 14.050 ;
        RECT 56.870 13.790 57.130 14.050 ;
        RECT 57.240 13.790 57.500 14.050 ;
        RECT 62.500 13.790 62.760 14.050 ;
        RECT 62.870 13.790 63.130 14.050 ;
        RECT 63.240 13.790 63.500 14.050 ;
        RECT 68.500 13.790 68.760 14.050 ;
        RECT 68.870 13.790 69.130 14.050 ;
        RECT 69.240 13.790 69.500 14.050 ;
        RECT 74.500 13.790 74.760 14.050 ;
        RECT 74.870 13.790 75.130 14.050 ;
        RECT 75.240 13.790 75.500 14.050 ;
        RECT 80.500 13.790 80.760 14.050 ;
        RECT 80.870 13.790 81.130 14.050 ;
        RECT 81.240 13.790 81.500 14.050 ;
        RECT 86.500 13.790 86.760 14.050 ;
        RECT 86.870 13.790 87.130 14.050 ;
        RECT 87.240 13.790 87.500 14.050 ;
        RECT 92.500 13.790 92.760 14.050 ;
        RECT 92.870 13.790 93.130 14.050 ;
        RECT 93.240 13.790 93.500 14.050 ;
        RECT 98.500 13.790 98.760 14.050 ;
        RECT 98.870 13.790 99.130 14.050 ;
        RECT 99.240 13.790 99.500 14.050 ;
        RECT 104.500 13.790 104.760 14.050 ;
        RECT 104.870 13.790 105.130 14.050 ;
        RECT 105.240 13.790 105.500 14.050 ;
        RECT 108.280 13.790 108.540 14.050 ;
        RECT 108.650 13.790 108.910 14.050 ;
        RECT 109.020 13.790 109.280 14.050 ;
      LAYER met2 ;
        RECT 104.500 18.500 105.500 19.515 ;
        RECT 14.500 15.700 15.500 16.100 ;
        RECT 20.500 15.700 21.500 16.100 ;
        RECT 26.500 15.700 27.500 16.100 ;
        RECT 32.500 15.700 33.500 16.100 ;
        RECT 38.500 15.700 39.500 16.100 ;
        RECT 44.500 15.700 45.500 16.100 ;
        RECT 50.500 15.700 51.500 16.100 ;
        RECT 56.500 15.700 57.500 16.100 ;
        RECT 62.500 15.700 63.500 16.100 ;
        RECT 68.500 15.700 69.500 16.100 ;
        RECT 74.500 15.700 75.500 16.100 ;
        RECT 80.500 15.700 81.500 16.100 ;
        RECT 86.500 15.700 87.500 16.100 ;
        RECT 92.500 15.700 93.500 16.100 ;
        RECT 98.500 15.700 99.500 16.100 ;
        RECT 2.500 13.720 3.500 14.120 ;
        RECT 8.500 13.720 9.500 14.120 ;
        RECT 14.500 13.720 15.500 14.120 ;
        RECT 20.500 13.720 21.500 14.120 ;
        RECT 26.500 13.720 27.500 14.120 ;
        RECT 32.500 13.720 33.500 14.120 ;
        RECT 38.500 13.720 39.500 14.120 ;
        RECT 44.500 13.720 45.500 14.120 ;
        RECT 50.500 13.720 51.500 14.120 ;
        RECT 56.500 13.720 57.500 14.120 ;
        RECT 62.500 13.720 63.500 14.120 ;
        RECT 68.500 13.720 69.500 14.120 ;
        RECT 74.500 13.720 75.500 14.120 ;
        RECT 80.500 13.720 81.500 14.120 ;
        RECT 86.500 13.720 87.500 14.120 ;
        RECT 92.500 13.720 93.500 14.120 ;
        RECT 98.500 13.720 99.500 14.120 ;
        RECT 104.500 13.720 105.500 14.120 ;
        RECT 108.280 13.720 109.280 14.120 ;
      LAYER via2 ;
        RECT 104.540 19.070 104.940 19.470 ;
        RECT 105.060 19.070 105.460 19.470 ;
        RECT 104.540 18.550 104.940 18.950 ;
        RECT 105.060 18.550 105.460 18.950 ;
        RECT 14.600 15.750 14.900 16.050 ;
        RECT 15.100 15.750 15.400 16.050 ;
        RECT 20.600 15.750 20.900 16.050 ;
        RECT 21.100 15.750 21.400 16.050 ;
        RECT 26.600 15.750 26.900 16.050 ;
        RECT 27.100 15.750 27.400 16.050 ;
        RECT 32.600 15.750 32.900 16.050 ;
        RECT 33.100 15.750 33.400 16.050 ;
        RECT 38.600 15.750 38.900 16.050 ;
        RECT 39.100 15.750 39.400 16.050 ;
        RECT 44.600 15.750 44.900 16.050 ;
        RECT 45.100 15.750 45.400 16.050 ;
        RECT 50.600 15.750 50.900 16.050 ;
        RECT 51.100 15.750 51.400 16.050 ;
        RECT 56.600 15.750 56.900 16.050 ;
        RECT 57.100 15.750 57.400 16.050 ;
        RECT 62.600 15.750 62.900 16.050 ;
        RECT 63.100 15.750 63.400 16.050 ;
        RECT 68.600 15.750 68.900 16.050 ;
        RECT 69.100 15.750 69.400 16.050 ;
        RECT 74.600 15.750 74.900 16.050 ;
        RECT 75.100 15.750 75.400 16.050 ;
        RECT 80.600 15.750 80.900 16.050 ;
        RECT 81.100 15.750 81.400 16.050 ;
        RECT 86.600 15.750 86.900 16.050 ;
        RECT 87.100 15.750 87.400 16.050 ;
        RECT 92.600 15.750 92.900 16.050 ;
        RECT 93.100 15.750 93.400 16.050 ;
        RECT 98.600 15.750 98.900 16.050 ;
        RECT 99.100 15.750 99.400 16.050 ;
        RECT 2.600 13.770 2.900 14.070 ;
        RECT 3.100 13.770 3.400 14.070 ;
        RECT 8.600 13.770 8.900 14.070 ;
        RECT 9.100 13.770 9.400 14.070 ;
        RECT 14.600 13.770 14.900 14.070 ;
        RECT 15.100 13.770 15.400 14.070 ;
        RECT 20.600 13.770 20.900 14.070 ;
        RECT 21.100 13.770 21.400 14.070 ;
        RECT 26.600 13.770 26.900 14.070 ;
        RECT 27.100 13.770 27.400 14.070 ;
        RECT 32.600 13.770 32.900 14.070 ;
        RECT 33.100 13.770 33.400 14.070 ;
        RECT 38.600 13.770 38.900 14.070 ;
        RECT 39.100 13.770 39.400 14.070 ;
        RECT 44.600 13.770 44.900 14.070 ;
        RECT 45.100 13.770 45.400 14.070 ;
        RECT 50.600 13.770 50.900 14.070 ;
        RECT 51.100 13.770 51.400 14.070 ;
        RECT 56.600 13.770 56.900 14.070 ;
        RECT 57.100 13.770 57.400 14.070 ;
        RECT 62.600 13.770 62.900 14.070 ;
        RECT 63.100 13.770 63.400 14.070 ;
        RECT 68.600 13.770 68.900 14.070 ;
        RECT 69.100 13.770 69.400 14.070 ;
        RECT 74.600 13.770 74.900 14.070 ;
        RECT 75.100 13.770 75.400 14.070 ;
        RECT 80.600 13.770 80.900 14.070 ;
        RECT 81.100 13.770 81.400 14.070 ;
        RECT 86.600 13.770 86.900 14.070 ;
        RECT 87.100 13.770 87.400 14.070 ;
        RECT 92.600 13.770 92.900 14.070 ;
        RECT 93.100 13.770 93.400 14.070 ;
        RECT 98.600 13.770 98.900 14.070 ;
        RECT 99.100 13.770 99.400 14.070 ;
        RECT 104.600 13.770 104.900 14.070 ;
        RECT 105.100 13.770 105.400 14.070 ;
        RECT 108.380 13.770 108.680 14.070 ;
        RECT 108.880 13.770 109.180 14.070 ;
      LAYER met3 ;
        RECT 14.500 15.670 15.500 16.150 ;
        RECT 20.500 15.670 21.500 16.150 ;
        RECT 26.500 15.670 27.500 16.150 ;
        RECT 32.500 15.670 33.500 16.150 ;
        RECT 38.500 15.670 39.500 16.150 ;
        RECT 44.500 15.670 45.500 16.150 ;
        RECT 50.500 15.670 51.500 16.150 ;
        RECT 56.500 15.670 57.500 16.150 ;
        RECT 62.500 15.670 63.500 16.150 ;
        RECT 68.500 15.670 69.500 16.150 ;
        RECT 74.500 15.670 75.500 16.150 ;
        RECT 80.500 15.670 81.500 16.150 ;
        RECT 86.500 15.670 87.500 16.150 ;
        RECT 92.500 15.670 93.500 16.150 ;
        RECT 98.500 15.670 99.500 16.150 ;
        RECT 104.500 15.670 105.500 19.515 ;
        RECT 2.500 14.170 109.280 15.670 ;
        RECT 2.500 13.690 3.500 14.170 ;
        RECT 8.500 13.690 9.500 14.170 ;
        RECT 14.500 13.690 15.500 14.170 ;
        RECT 20.500 13.690 21.500 14.170 ;
        RECT 26.500 13.690 27.500 14.170 ;
        RECT 32.500 13.690 33.500 14.170 ;
        RECT 38.500 13.690 39.500 14.170 ;
        RECT 44.500 13.690 45.500 14.170 ;
        RECT 50.500 13.690 51.500 14.170 ;
        RECT 56.500 13.690 57.500 14.170 ;
        RECT 62.500 13.690 63.500 14.170 ;
        RECT 68.500 13.690 69.500 14.170 ;
        RECT 74.500 13.690 75.500 14.170 ;
        RECT 80.500 13.690 81.500 14.170 ;
        RECT 86.500 13.690 87.500 14.170 ;
        RECT 92.500 13.690 93.500 14.170 ;
        RECT 98.500 13.690 99.500 14.170 ;
        RECT 104.500 13.690 105.500 14.170 ;
        RECT 108.280 13.690 109.280 14.170 ;
  END
END vco_w6_r100
END LIBRARY

