magic
tech sky130A
magscale 1 2
timestamp 1637949574
<< pwell >>
rect 1601 12232 1687 12318
<< ndiff >>
rect 1627 12258 1661 12292
<< pdiff >>
rect 1627 12582 1661 12616
<< locali >>
rect 1910 12548 1955 12592
rect 2308 12542 2353 12586
rect 600 12467 1356 12480
rect 600 12433 613 12467
rect 647 12433 1356 12467
rect 600 12420 1356 12433
rect 1496 12384 1521 12418
<< viali >>
rect 613 12433 647 12467
<< metal1 >>
rect 0 12656 1994 12752
rect 598 12476 662 12482
rect 598 12424 604 12476
rect 656 12424 662 12476
rect 598 12418 662 12424
rect 5898 12452 5970 12462
rect 5898 12400 5908 12452
rect 5960 12400 5970 12452
rect 5898 12390 5970 12400
rect 10568 12452 10652 12462
rect 10568 12400 10584 12452
rect 10636 12400 10652 12452
rect 10568 12390 10652 12400
rect 14110 12452 14194 12462
rect 14110 12400 14126 12452
rect 14178 12400 14194 12452
rect 14110 12390 14194 12400
rect 16656 12452 16740 12462
rect 16656 12400 16672 12452
rect 16724 12400 16740 12452
rect 16656 12390 16740 12400
rect 21082 12452 21382 12462
rect 21082 12400 21180 12452
rect 21232 12400 21382 12452
rect 21722 12404 23600 12476
rect 21082 12390 21382 12400
rect 800 12112 1962 12208
rect 1226 8768 1562 8778
rect 1226 8716 1400 8768
rect 1452 8716 1562 8768
rect 1226 8706 1562 8716
rect 4774 8768 4858 8778
rect 4774 8716 4790 8768
rect 4842 8716 4858 8768
rect 4774 8706 4858 8716
rect 8560 8768 8644 8778
rect 8560 8716 8576 8768
rect 8628 8716 8644 8768
rect 8560 8706 8644 8716
rect 13160 8768 13244 8778
rect 13160 8716 13176 8768
rect 13228 8716 13244 8768
rect 13160 8706 13244 8716
rect 15644 8768 15728 8778
rect 15644 8716 15660 8768
rect 15712 8716 15728 8768
rect 15644 8706 15728 8716
rect 19232 8768 19316 8778
rect 19232 8716 19248 8768
rect 19300 8716 19316 8768
rect 19232 8706 19316 8716
<< via1 >>
rect 604 12467 656 12476
rect 604 12433 613 12467
rect 613 12433 647 12467
rect 647 12433 656 12467
rect 604 12424 656 12433
rect 5908 12400 5960 12452
rect 10584 12400 10636 12452
rect 14126 12400 14178 12452
rect 16672 12400 16724 12452
rect 21180 12400 21232 12452
rect 1400 8716 1452 8768
rect 4790 8716 4842 8768
rect 8576 8716 8628 8768
rect 13176 8716 13228 8768
rect 15660 8716 15712 8768
rect 19248 8716 19300 8768
<< metal2 >>
rect 590 12478 670 12480
rect 590 12422 602 12478
rect 658 12422 670 12478
rect 590 12420 670 12422
rect 5842 12452 6026 12472
rect 5842 12400 5908 12452
rect 5960 12400 6026 12452
rect 5842 12380 6026 12400
rect 10518 12452 10702 12472
rect 10518 12400 10584 12452
rect 10636 12400 10702 12452
rect 10518 12380 10702 12400
rect 14060 12452 14244 12472
rect 14060 12400 14126 12452
rect 14178 12400 14244 12452
rect 14060 12380 14244 12400
rect 16606 12452 16790 12472
rect 16606 12400 16672 12452
rect 16724 12400 16790 12452
rect 16606 12380 16790 12400
rect 21114 12452 21298 12472
rect 21114 12400 21180 12452
rect 21232 12400 21298 12452
rect 21114 12380 21298 12400
rect 24426 11520 24610 11542
rect 24426 11464 24490 11520
rect 24546 11464 24610 11520
rect 24426 11442 24610 11464
rect 1334 8768 1518 8788
rect 1334 8716 1400 8768
rect 1452 8716 1518 8768
rect 1334 8696 1518 8716
rect 4724 8768 4908 8788
rect 4724 8716 4790 8768
rect 4842 8716 4908 8768
rect 4724 8696 4908 8716
rect 8510 8768 8694 8788
rect 8510 8716 8576 8768
rect 8628 8716 8694 8768
rect 8510 8696 8694 8716
rect 13110 8768 13294 8788
rect 13110 8716 13176 8768
rect 13228 8716 13294 8768
rect 13110 8696 13294 8716
rect 15594 8768 15778 8788
rect 15594 8716 15660 8768
rect 15712 8716 15778 8768
rect 15594 8696 15778 8716
rect 19182 8768 19366 8788
rect 19182 8716 19248 8768
rect 19300 8716 19366 8768
rect 19182 8696 19366 8716
<< via2 >>
rect 602 12476 658 12478
rect 602 12424 604 12476
rect 604 12424 656 12476
rect 656 12424 658 12476
rect 602 12422 658 12424
rect 24490 11464 24546 11520
<< metal3 >>
rect 0 20600 5200 21000
rect 590 12930 670 13010
rect 592 12478 668 12930
rect 592 12422 602 12478
rect 658 12422 668 12478
rect 592 12412 668 12422
rect 24464 11520 24572 11628
rect 24464 11464 24490 11520
rect 24546 11464 24572 11520
rect 24464 11356 24572 11464
rect 18600 800 23600 1200
use pwell_co_ring_w6  pwell_co_ring_w6_0
timestamp 1623529308
transform 1 0 3020 0 1 13740
box -1680 -6360 20145 60
use via_m4_li  via_m4_li_0
timestamp 1623563441
transform 1 0 12000 0 1 7360
box 0 2 400 98
use via_m4_li  via_m4_li_1
timestamp 1623563441
transform 1 0 6400 0 1 7360
box 0 2 400 98
use via_m1  via_m1_0
timestamp 1623561200
transform 1 0 9502 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_1
timestamp 1623561200
transform 1 0 3902 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_2
timestamp 1623561200
transform 1 0 -1698 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_3
timestamp 1623561200
transform 1 0 -7298 0 1 662
box 10898 6956 11298 7052
use ring_osc_w6  ring_osc_w6_0
timestamp 1637949574
transform 1 0 1500 0 1 7600
box -502 0 23110 5968
use via_m1  via_m1_4
timestamp 1623561200
transform 1 0 -10898 0 1 5700
box 10898 6956 11298 7052
use via_m1  via_m1_5
timestamp 1623561200
transform 1 0 -10098 0 1 5156
box 10898 6956 11298 7052
use via_m1  via_m1_6
timestamp 1623561200
transform 1 0 -7298 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_2
timestamp 1623563441
transform 1 0 6400 0 1 13720
box 0 2 400 98
use via_m1  via_m1_7
timestamp 1623561200
transform 1 0 -1698 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_3
timestamp 1623563441
transform 1 0 12000 0 1 13720
box 0 2 400 98
use via_m1  via_m1_8
timestamp 1623561200
transform 1 0 3902 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_4
timestamp 1623563441
transform 1 0 17600 0 1 13720
box 0 2 400 98
use via_m1  via_m1_9
timestamp 1623561200
transform 1 0 12302 0 1 5436
box 10898 6956 11298 7052
use via_m1  via_m1_10
timestamp 1623561200
transform 1 0 9502 0 1 6498
box 10898 6956 11298 7052
use power_ring  power_ring_0
timestamp 1623530672
transform 1 0 0 0 1 0
box 0 0 24400 21000
<< labels >>
flabel metal2 s 19232 8700 19316 8784 1 FreeSans 800 0 0 0 p[9]
port 1 nsew signal output
flabel metal2 s 15644 8700 15728 8784 1 FreeSans 800 0 0 0 p[7]
port 2 nsew signal output
flabel metal2 s 13160 8700 13244 8784 1 FreeSans 800 0 0 0 p[5]
port 3 nsew signal output
flabel metal2 s 8560 8700 8644 8784 1 FreeSans 800 0 0 0 p[3]
port 4 nsew signal output
flabel metal2 s 4774 8700 4858 8784 1 FreeSans 800 0 0 0 p[1]
port 5 nsew signal output
flabel metal2 s 1384 8700 1468 8784 1 FreeSans 800 0 0 0 p[0]
port 6 nsew signal output
flabel metal2 s 5892 12384 5976 12468 1 FreeSans 800 0 0 0 p[2]
port 7 nsew signal output
flabel metal2 s 10568 12384 10652 12468 1 FreeSans 800 0 0 0 p[4]
port 8 nsew signal output
flabel metal2 s 14110 12384 14194 12468 1 FreeSans 800 0 0 0 p[6]
port 9 nsew signal output
flabel metal2 s 16656 12384 16740 12468 1 FreeSans 800 0 0 0 p[8]
port 10 nsew signal output
flabel metal2 s 21164 12384 21248 12468 1 FreeSans 800 0 0 0 p[10]
port 11 nsew signal output
flabel metal3 s 590 12930 670 13010 1 FreeSans 800 0 0 0 enb
port 12 nsew signal input
flabel metal2 s 24468 11442 24568 11542 1 FreeSans 800 0 0 0 input_analog
port 13 nsew signal input
flabel metal3 s 0 20600 5200 21000 1 FreeSans 20 0 0 0 vccd2
port 14 nsew power bidirectional 
flabel metal3 s 18600 800 23600 1200 1 FreeSans 20 0 0 0 vssd2
port 15 nsew ground bidirectional
<< end >>
