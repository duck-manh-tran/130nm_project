magic
tech sky130A
magscale 1 2
timestamp 1623147637
<< nwell >>
rect 0 -2 772 1374
<< pmos >>
rect 196 217 576 1217
<< pdiff >>
rect 138 1181 196 1217
rect 138 1141 150 1181
rect 184 1141 196 1181
rect 138 1107 196 1141
rect 138 1067 150 1107
rect 184 1067 196 1107
rect 138 1033 196 1067
rect 138 993 150 1033
rect 184 993 196 1033
rect 138 959 196 993
rect 138 919 150 959
rect 184 919 196 959
rect 138 885 196 919
rect 138 845 150 885
rect 184 845 196 885
rect 138 811 196 845
rect 138 771 150 811
rect 184 771 196 811
rect 138 737 196 771
rect 138 697 150 737
rect 184 697 196 737
rect 138 663 196 697
rect 138 623 150 663
rect 184 623 196 663
rect 138 589 196 623
rect 138 549 150 589
rect 184 549 196 589
rect 138 515 196 549
rect 138 475 150 515
rect 184 475 196 515
rect 138 441 196 475
rect 138 401 150 441
rect 184 401 196 441
rect 138 367 196 401
rect 138 327 150 367
rect 184 327 196 367
rect 138 293 196 327
rect 138 253 150 293
rect 184 253 196 293
rect 138 217 196 253
rect 576 1181 634 1217
rect 576 1141 588 1181
rect 622 1141 634 1181
rect 576 1107 634 1141
rect 576 1067 588 1107
rect 622 1067 634 1107
rect 576 1033 634 1067
rect 576 993 588 1033
rect 622 993 634 1033
rect 576 959 634 993
rect 576 919 588 959
rect 622 919 634 959
rect 576 885 634 919
rect 576 845 588 885
rect 622 845 634 885
rect 576 811 634 845
rect 576 771 588 811
rect 622 771 634 811
rect 576 737 634 771
rect 576 697 588 737
rect 622 697 634 737
rect 576 663 634 697
rect 576 623 588 663
rect 622 623 634 663
rect 576 589 634 623
rect 576 549 588 589
rect 622 549 634 589
rect 576 515 634 549
rect 576 475 588 515
rect 622 475 634 515
rect 576 441 634 475
rect 576 401 588 441
rect 622 401 634 441
rect 576 367 634 401
rect 576 327 588 367
rect 622 327 634 367
rect 576 293 634 327
rect 576 253 588 293
rect 622 253 634 293
rect 576 217 634 253
<< pdiffc >>
rect 150 1141 184 1181
rect 150 1067 184 1107
rect 150 993 184 1033
rect 150 919 184 959
rect 150 845 184 885
rect 150 771 184 811
rect 150 697 184 737
rect 150 623 184 663
rect 150 549 184 589
rect 150 475 184 515
rect 150 401 184 441
rect 150 327 184 367
rect 150 253 184 293
rect 588 1141 622 1181
rect 588 1067 622 1107
rect 588 993 622 1033
rect 588 919 622 959
rect 588 845 622 885
rect 588 771 622 811
rect 588 697 622 737
rect 588 623 622 663
rect 588 549 622 589
rect 588 475 622 515
rect 588 401 622 441
rect 588 327 622 367
rect 588 253 622 293
<< nsubdiff >>
rect 36 1304 140 1338
rect 180 1304 220 1338
rect 260 1304 300 1338
rect 340 1304 380 1338
rect 420 1304 460 1338
rect 500 1304 540 1338
rect 580 1304 620 1338
rect 660 1304 736 1338
<< nsubdiffcont >>
rect 140 1304 180 1338
rect 220 1304 260 1338
rect 300 1304 340 1338
rect 380 1304 420 1338
rect 460 1304 500 1338
rect 540 1304 580 1338
rect 620 1304 660 1338
<< poly >>
rect 196 1217 576 1243
rect 196 120 576 217
<< locali >>
rect 36 1304 140 1338
rect 180 1304 220 1338
rect 260 1304 300 1338
rect 340 1304 380 1338
rect 420 1304 460 1338
rect 500 1304 540 1338
rect 580 1304 620 1338
rect 660 1304 736 1338
rect 138 1181 196 1304
rect 138 1141 150 1181
rect 184 1141 196 1181
rect 138 1107 196 1141
rect 138 1067 150 1107
rect 184 1067 196 1107
rect 138 1033 196 1067
rect 138 993 150 1033
rect 184 993 196 1033
rect 138 959 196 993
rect 138 919 150 959
rect 184 919 196 959
rect 138 885 196 919
rect 138 845 150 885
rect 184 845 196 885
rect 138 811 196 845
rect 138 771 150 811
rect 184 771 196 811
rect 138 737 196 771
rect 138 697 150 737
rect 184 697 196 737
rect 138 663 196 697
rect 138 623 150 663
rect 184 623 196 663
rect 138 589 196 623
rect 138 549 150 589
rect 184 549 196 589
rect 138 515 196 549
rect 138 475 150 515
rect 184 475 196 515
rect 138 441 196 475
rect 138 401 150 441
rect 184 401 196 441
rect 138 367 196 401
rect 138 327 150 367
rect 184 327 196 367
rect 138 293 196 327
rect 138 253 150 293
rect 184 253 196 293
rect 138 212 196 253
rect 588 1181 622 1221
rect 588 1107 622 1141
rect 588 1033 622 1067
rect 588 959 622 993
rect 588 885 622 919
rect 588 811 622 845
rect 588 737 622 771
rect 588 663 622 697
rect 588 589 622 623
rect 588 515 622 549
rect 588 441 622 475
rect 588 367 622 401
rect 588 293 622 327
rect 588 213 622 253
<< end >>
