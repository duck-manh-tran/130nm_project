magic
tech sky130A
timestamp 1623991673
<< metal3 >>
rect 15300 12080 29880 12100
rect 15300 12040 15320 12080
rect 15360 12040 15380 12080
rect 15420 12040 15440 12080
rect 15480 12040 18920 12080
rect 18960 12040 18980 12080
rect 19020 12040 19040 12080
rect 19080 12040 22520 12080
rect 22560 12040 22580 12080
rect 22620 12040 22640 12080
rect 22680 12040 26120 12080
rect 26160 12040 26180 12080
rect 26220 12040 26240 12080
rect 26280 12040 29720 12080
rect 29760 12040 29780 12080
rect 29820 12040 29840 12080
rect 15300 12020 29880 12040
rect 15300 11980 15320 12020
rect 15360 11980 15380 12020
rect 15420 11980 15440 12020
rect 15480 11980 18920 12020
rect 18960 11980 18980 12020
rect 19020 11980 19040 12020
rect 19080 11980 22520 12020
rect 22560 11980 22580 12020
rect 22620 11980 22640 12020
rect 22680 11980 26120 12020
rect 26160 11980 26180 12020
rect 26220 11980 26240 12020
rect 26280 11980 29720 12020
rect 29760 11980 29780 12020
rect 29820 11980 29840 12020
rect 15300 11960 29880 11980
rect 15300 11920 15320 11960
rect 15360 11920 15380 11960
rect 15420 11920 15440 11960
rect 15480 11920 18920 11960
rect 18960 11920 18980 11960
rect 19020 11920 19040 11960
rect 19080 11920 22520 11960
rect 22560 11920 22580 11960
rect 22620 11920 22640 11960
rect 22680 11920 26120 11960
rect 26160 11920 26180 11960
rect 26220 11920 26240 11960
rect 26280 11920 29720 11960
rect 29760 11920 29780 11960
rect 29820 11920 29840 11960
rect 15300 11900 29880 11920
rect 13500 11680 31700 11700
rect 13500 11640 13520 11680
rect 13560 11640 13580 11680
rect 13620 11640 13640 11680
rect 13680 11640 17120 11680
rect 17160 11640 17180 11680
rect 17220 11640 17240 11680
rect 17280 11640 20720 11680
rect 20760 11640 20780 11680
rect 20820 11640 20840 11680
rect 20880 11640 24320 11680
rect 24360 11640 24380 11680
rect 24420 11640 24440 11680
rect 24480 11640 27920 11680
rect 27960 11640 27980 11680
rect 28020 11640 28040 11680
rect 28080 11640 31520 11680
rect 31560 11640 31580 11680
rect 31620 11640 31640 11680
rect 31680 11640 31700 11680
rect 13500 11620 31700 11640
rect 13500 11580 13520 11620
rect 13560 11580 13580 11620
rect 13620 11580 13640 11620
rect 13680 11580 17120 11620
rect 17160 11580 17180 11620
rect 17220 11580 17240 11620
rect 17280 11580 20720 11620
rect 20760 11580 20780 11620
rect 20820 11580 20840 11620
rect 20880 11580 24320 11620
rect 24360 11580 24380 11620
rect 24420 11580 24440 11620
rect 24480 11580 27920 11620
rect 27960 11580 27980 11620
rect 28020 11580 28040 11620
rect 28080 11580 31520 11620
rect 31560 11580 31580 11620
rect 31620 11580 31640 11620
rect 31680 11580 31700 11620
rect 13500 11560 31700 11580
rect 13500 11520 13520 11560
rect 13560 11520 13580 11560
rect 13620 11520 13640 11560
rect 13680 11520 17120 11560
rect 17160 11520 17180 11560
rect 17220 11520 17240 11560
rect 17280 11520 20720 11560
rect 20760 11520 20780 11560
rect 20820 11520 20840 11560
rect 20880 11520 24320 11560
rect 24360 11520 24380 11560
rect 24420 11520 24440 11560
rect 24480 11520 27920 11560
rect 27960 11520 27980 11560
rect 28020 11520 28040 11560
rect 28080 11520 31520 11560
rect 31560 11520 31580 11560
rect 31620 11520 31640 11560
rect 31680 11520 31700 11560
rect 13500 11500 31700 11520
rect 13500 2180 31700 2200
rect 13500 2140 13520 2180
rect 13560 2140 13580 2180
rect 13620 2140 13640 2180
rect 13680 2140 17120 2180
rect 17160 2140 17180 2180
rect 17220 2140 17240 2180
rect 17280 2140 20720 2180
rect 20760 2140 20780 2180
rect 20820 2140 20840 2180
rect 20880 2140 24320 2180
rect 24360 2140 24380 2180
rect 24420 2140 24440 2180
rect 24480 2140 27920 2180
rect 27960 2140 27980 2180
rect 28020 2140 28040 2180
rect 28080 2140 31520 2180
rect 31560 2140 31580 2180
rect 31620 2140 31640 2180
rect 31680 2140 31700 2180
rect 13500 2120 31700 2140
rect 13500 2080 13520 2120
rect 13560 2080 13580 2120
rect 13620 2080 13640 2120
rect 13680 2080 17120 2120
rect 17160 2080 17180 2120
rect 17220 2080 17240 2120
rect 17280 2080 20720 2120
rect 20760 2080 20780 2120
rect 20820 2080 20840 2120
rect 20880 2080 24320 2120
rect 24360 2080 24380 2120
rect 24420 2080 24440 2120
rect 24480 2080 27920 2120
rect 27960 2080 27980 2120
rect 28020 2080 28040 2120
rect 28080 2080 31520 2120
rect 31560 2080 31580 2120
rect 31620 2080 31640 2120
rect 31680 2080 31700 2120
rect 13500 2060 31700 2080
rect 13500 2020 13520 2060
rect 13560 2020 13580 2060
rect 13620 2020 13640 2060
rect 13680 2020 17120 2060
rect 17160 2020 17180 2060
rect 17220 2020 17240 2060
rect 17280 2020 20720 2060
rect 20760 2020 20780 2060
rect 20820 2020 20840 2060
rect 20880 2020 24320 2060
rect 24360 2020 24380 2060
rect 24420 2020 24440 2060
rect 24480 2020 27920 2060
rect 27960 2020 27980 2060
rect 28020 2020 28040 2060
rect 28080 2020 31520 2060
rect 31560 2020 31580 2060
rect 31620 2020 31640 2060
rect 31680 2020 31700 2060
rect 13500 2000 31700 2020
rect 15300 1780 29880 1800
rect 15300 1740 15320 1780
rect 15360 1740 15380 1780
rect 15420 1740 15440 1780
rect 15480 1740 18920 1780
rect 18960 1740 18980 1780
rect 19020 1740 19040 1780
rect 19080 1740 22520 1780
rect 22560 1740 22580 1780
rect 22620 1740 22640 1780
rect 22680 1740 26120 1780
rect 26160 1740 26180 1780
rect 26220 1740 26240 1780
rect 26280 1740 29720 1780
rect 29760 1740 29780 1780
rect 29820 1740 29840 1780
rect 15300 1720 29880 1740
rect 15300 1680 15320 1720
rect 15360 1680 15380 1720
rect 15420 1680 15440 1720
rect 15480 1680 18920 1720
rect 18960 1680 18980 1720
rect 19020 1680 19040 1720
rect 19080 1680 22520 1720
rect 22560 1680 22580 1720
rect 22620 1680 22640 1720
rect 22680 1680 26120 1720
rect 26160 1680 26180 1720
rect 26220 1680 26240 1720
rect 26280 1680 29720 1720
rect 29760 1680 29780 1720
rect 29820 1680 29840 1720
rect 15300 1660 29880 1680
rect 15300 1620 15320 1660
rect 15360 1620 15380 1660
rect 15420 1620 15440 1660
rect 15480 1620 18920 1660
rect 18960 1620 18980 1660
rect 19020 1620 19040 1660
rect 19080 1620 22520 1660
rect 22560 1620 22580 1660
rect 22620 1620 22640 1660
rect 22680 1620 26120 1660
rect 26160 1620 26180 1660
rect 26220 1620 26240 1660
rect 26280 1620 29720 1660
rect 29760 1620 29780 1660
rect 29820 1620 29840 1660
rect 15300 1600 29880 1620
<< via3 >>
rect 15320 12040 15360 12080
rect 15380 12040 15420 12080
rect 15440 12040 15480 12080
rect 18920 12040 18960 12080
rect 18980 12040 19020 12080
rect 19040 12040 19080 12080
rect 22520 12040 22560 12080
rect 22580 12040 22620 12080
rect 22640 12040 22680 12080
rect 26120 12040 26160 12080
rect 26180 12040 26220 12080
rect 26240 12040 26280 12080
rect 29720 12040 29760 12080
rect 29780 12040 29820 12080
rect 29840 12040 29880 12080
rect 15320 11980 15360 12020
rect 15380 11980 15420 12020
rect 15440 11980 15480 12020
rect 18920 11980 18960 12020
rect 18980 11980 19020 12020
rect 19040 11980 19080 12020
rect 22520 11980 22560 12020
rect 22580 11980 22620 12020
rect 22640 11980 22680 12020
rect 26120 11980 26160 12020
rect 26180 11980 26220 12020
rect 26240 11980 26280 12020
rect 29720 11980 29760 12020
rect 29780 11980 29820 12020
rect 29840 11980 29880 12020
rect 15320 11920 15360 11960
rect 15380 11920 15420 11960
rect 15440 11920 15480 11960
rect 18920 11920 18960 11960
rect 18980 11920 19020 11960
rect 19040 11920 19080 11960
rect 22520 11920 22560 11960
rect 22580 11920 22620 11960
rect 22640 11920 22680 11960
rect 26120 11920 26160 11960
rect 26180 11920 26220 11960
rect 26240 11920 26280 11960
rect 29720 11920 29760 11960
rect 29780 11920 29820 11960
rect 29840 11920 29880 11960
rect 13520 11640 13560 11680
rect 13580 11640 13620 11680
rect 13640 11640 13680 11680
rect 17120 11640 17160 11680
rect 17180 11640 17220 11680
rect 17240 11640 17280 11680
rect 20720 11640 20760 11680
rect 20780 11640 20820 11680
rect 20840 11640 20880 11680
rect 24320 11640 24360 11680
rect 24380 11640 24420 11680
rect 24440 11640 24480 11680
rect 27920 11640 27960 11680
rect 27980 11640 28020 11680
rect 28040 11640 28080 11680
rect 31520 11640 31560 11680
rect 31580 11640 31620 11680
rect 31640 11640 31680 11680
rect 13520 11580 13560 11620
rect 13580 11580 13620 11620
rect 13640 11580 13680 11620
rect 17120 11580 17160 11620
rect 17180 11580 17220 11620
rect 17240 11580 17280 11620
rect 20720 11580 20760 11620
rect 20780 11580 20820 11620
rect 20840 11580 20880 11620
rect 24320 11580 24360 11620
rect 24380 11580 24420 11620
rect 24440 11580 24480 11620
rect 27920 11580 27960 11620
rect 27980 11580 28020 11620
rect 28040 11580 28080 11620
rect 31520 11580 31560 11620
rect 31580 11580 31620 11620
rect 31640 11580 31680 11620
rect 13520 11520 13560 11560
rect 13580 11520 13620 11560
rect 13640 11520 13680 11560
rect 17120 11520 17160 11560
rect 17180 11520 17220 11560
rect 17240 11520 17280 11560
rect 20720 11520 20760 11560
rect 20780 11520 20820 11560
rect 20840 11520 20880 11560
rect 24320 11520 24360 11560
rect 24380 11520 24420 11560
rect 24440 11520 24480 11560
rect 27920 11520 27960 11560
rect 27980 11520 28020 11560
rect 28040 11520 28080 11560
rect 31520 11520 31560 11560
rect 31580 11520 31620 11560
rect 31640 11520 31680 11560
rect 13520 2140 13560 2180
rect 13580 2140 13620 2180
rect 13640 2140 13680 2180
rect 17120 2140 17160 2180
rect 17180 2140 17220 2180
rect 17240 2140 17280 2180
rect 20720 2140 20760 2180
rect 20780 2140 20820 2180
rect 20840 2140 20880 2180
rect 24320 2140 24360 2180
rect 24380 2140 24420 2180
rect 24440 2140 24480 2180
rect 27920 2140 27960 2180
rect 27980 2140 28020 2180
rect 28040 2140 28080 2180
rect 31520 2140 31560 2180
rect 31580 2140 31620 2180
rect 31640 2140 31680 2180
rect 13520 2080 13560 2120
rect 13580 2080 13620 2120
rect 13640 2080 13680 2120
rect 17120 2080 17160 2120
rect 17180 2080 17220 2120
rect 17240 2080 17280 2120
rect 20720 2080 20760 2120
rect 20780 2080 20820 2120
rect 20840 2080 20880 2120
rect 24320 2080 24360 2120
rect 24380 2080 24420 2120
rect 24440 2080 24480 2120
rect 27920 2080 27960 2120
rect 27980 2080 28020 2120
rect 28040 2080 28080 2120
rect 31520 2080 31560 2120
rect 31580 2080 31620 2120
rect 31640 2080 31680 2120
rect 13520 2020 13560 2060
rect 13580 2020 13620 2060
rect 13640 2020 13680 2060
rect 17120 2020 17160 2060
rect 17180 2020 17220 2060
rect 17240 2020 17280 2060
rect 20720 2020 20760 2060
rect 20780 2020 20820 2060
rect 20840 2020 20880 2060
rect 24320 2020 24360 2060
rect 24380 2020 24420 2060
rect 24440 2020 24480 2060
rect 27920 2020 27960 2060
rect 27980 2020 28020 2060
rect 28040 2020 28080 2060
rect 31520 2020 31560 2060
rect 31580 2020 31620 2060
rect 31640 2020 31680 2060
rect 15320 1740 15360 1780
rect 15380 1740 15420 1780
rect 15440 1740 15480 1780
rect 18920 1740 18960 1780
rect 18980 1740 19020 1780
rect 19040 1740 19080 1780
rect 22520 1740 22560 1780
rect 22580 1740 22620 1780
rect 22640 1740 22680 1780
rect 26120 1740 26160 1780
rect 26180 1740 26220 1780
rect 26240 1740 26280 1780
rect 29720 1740 29760 1780
rect 29780 1740 29820 1780
rect 29840 1740 29880 1780
rect 15320 1680 15360 1720
rect 15380 1680 15420 1720
rect 15440 1680 15480 1720
rect 18920 1680 18960 1720
rect 18980 1680 19020 1720
rect 19040 1680 19080 1720
rect 22520 1680 22560 1720
rect 22580 1680 22620 1720
rect 22640 1680 22680 1720
rect 26120 1680 26160 1720
rect 26180 1680 26220 1720
rect 26240 1680 26280 1720
rect 29720 1680 29760 1720
rect 29780 1680 29820 1720
rect 29840 1680 29880 1720
rect 15320 1620 15360 1660
rect 15380 1620 15420 1660
rect 15440 1620 15480 1660
rect 18920 1620 18960 1660
rect 18980 1620 19020 1660
rect 19040 1620 19080 1660
rect 22520 1620 22560 1660
rect 22580 1620 22620 1660
rect 22640 1620 22680 1660
rect 26120 1620 26160 1660
rect 26180 1620 26220 1660
rect 26240 1620 26280 1660
rect 29720 1620 29760 1660
rect 29780 1620 29820 1660
rect 29840 1620 29880 1660
<< metal4 >>
rect 15300 12080 15500 12100
rect 15300 12040 15320 12080
rect 15360 12040 15380 12080
rect 15420 12040 15440 12080
rect 15480 12040 15500 12080
rect 15300 12020 15500 12040
rect 15300 11980 15320 12020
rect 15360 11980 15380 12020
rect 15420 11980 15440 12020
rect 15480 11980 15500 12020
rect 15300 11960 15500 11980
rect 15300 11920 15320 11960
rect 15360 11920 15380 11960
rect 15420 11920 15440 11960
rect 15480 11920 15500 11960
rect 13500 11680 13700 11700
rect 13500 11640 13520 11680
rect 13560 11640 13580 11680
rect 13620 11640 13640 11680
rect 13680 11640 13700 11680
rect 13500 11620 13700 11640
rect 13500 11580 13520 11620
rect 13560 11580 13580 11620
rect 13620 11580 13640 11620
rect 13680 11580 13700 11620
rect 13500 11560 13700 11580
rect 13500 11520 13520 11560
rect 13560 11520 13580 11560
rect 13620 11520 13640 11560
rect 13680 11520 13700 11560
rect 13500 2180 13700 11520
rect 13500 2140 13520 2180
rect 13560 2140 13580 2180
rect 13620 2140 13640 2180
rect 13680 2140 13700 2180
rect 13500 2120 13700 2140
rect 13500 2080 13520 2120
rect 13560 2080 13580 2120
rect 13620 2080 13640 2120
rect 13680 2080 13700 2120
rect 13500 2060 13700 2080
rect 13500 2020 13520 2060
rect 13560 2020 13580 2060
rect 13620 2020 13640 2060
rect 13680 2020 13700 2060
rect 13500 2000 13700 2020
rect 15300 1780 15500 11920
rect 18900 12080 19100 12100
rect 18900 12040 18920 12080
rect 18960 12040 18980 12080
rect 19020 12040 19040 12080
rect 19080 12040 19100 12080
rect 18900 12020 19100 12040
rect 18900 11980 18920 12020
rect 18960 11980 18980 12020
rect 19020 11980 19040 12020
rect 19080 11980 19100 12020
rect 18900 11960 19100 11980
rect 18900 11920 18920 11960
rect 18960 11920 18980 11960
rect 19020 11920 19040 11960
rect 19080 11920 19100 11960
rect 17100 11680 17300 11700
rect 17100 11640 17120 11680
rect 17160 11640 17180 11680
rect 17220 11640 17240 11680
rect 17280 11640 17300 11680
rect 17100 11620 17300 11640
rect 17100 11580 17120 11620
rect 17160 11580 17180 11620
rect 17220 11580 17240 11620
rect 17280 11580 17300 11620
rect 17100 11560 17300 11580
rect 17100 11520 17120 11560
rect 17160 11520 17180 11560
rect 17220 11520 17240 11560
rect 17280 11520 17300 11560
rect 17100 2180 17300 11520
rect 17100 2140 17120 2180
rect 17160 2140 17180 2180
rect 17220 2140 17240 2180
rect 17280 2140 17300 2180
rect 17100 2120 17300 2140
rect 17100 2080 17120 2120
rect 17160 2080 17180 2120
rect 17220 2080 17240 2120
rect 17280 2080 17300 2120
rect 17100 2060 17300 2080
rect 17100 2020 17120 2060
rect 17160 2020 17180 2060
rect 17220 2020 17240 2060
rect 17280 2020 17300 2060
rect 17100 2000 17300 2020
rect 15300 1740 15320 1780
rect 15360 1740 15380 1780
rect 15420 1740 15440 1780
rect 15480 1740 15500 1780
rect 15300 1720 15500 1740
rect 15300 1680 15320 1720
rect 15360 1680 15380 1720
rect 15420 1680 15440 1720
rect 15480 1680 15500 1720
rect 15300 1660 15500 1680
rect 15300 1620 15320 1660
rect 15360 1620 15380 1660
rect 15420 1620 15440 1660
rect 15480 1620 15500 1660
rect 15300 1600 15500 1620
rect 18900 1780 19100 11920
rect 22500 12080 22700 12100
rect 22500 12040 22520 12080
rect 22560 12040 22580 12080
rect 22620 12040 22640 12080
rect 22680 12040 22700 12080
rect 22500 12020 22700 12040
rect 22500 11980 22520 12020
rect 22560 11980 22580 12020
rect 22620 11980 22640 12020
rect 22680 11980 22700 12020
rect 22500 11960 22700 11980
rect 22500 11920 22520 11960
rect 22560 11920 22580 11960
rect 22620 11920 22640 11960
rect 22680 11920 22700 11960
rect 20700 11680 20900 11700
rect 20700 11640 20720 11680
rect 20760 11640 20780 11680
rect 20820 11640 20840 11680
rect 20880 11640 20900 11680
rect 20700 11620 20900 11640
rect 20700 11580 20720 11620
rect 20760 11580 20780 11620
rect 20820 11580 20840 11620
rect 20880 11580 20900 11620
rect 20700 11560 20900 11580
rect 20700 11520 20720 11560
rect 20760 11520 20780 11560
rect 20820 11520 20840 11560
rect 20880 11520 20900 11560
rect 20700 2180 20900 11520
rect 20700 2140 20720 2180
rect 20760 2140 20780 2180
rect 20820 2140 20840 2180
rect 20880 2140 20900 2180
rect 20700 2120 20900 2140
rect 20700 2080 20720 2120
rect 20760 2080 20780 2120
rect 20820 2080 20840 2120
rect 20880 2080 20900 2120
rect 20700 2060 20900 2080
rect 20700 2020 20720 2060
rect 20760 2020 20780 2060
rect 20820 2020 20840 2060
rect 20880 2020 20900 2060
rect 20700 2000 20900 2020
rect 18900 1740 18920 1780
rect 18960 1740 18980 1780
rect 19020 1740 19040 1780
rect 19080 1740 19100 1780
rect 18900 1720 19100 1740
rect 18900 1680 18920 1720
rect 18960 1680 18980 1720
rect 19020 1680 19040 1720
rect 19080 1680 19100 1720
rect 18900 1660 19100 1680
rect 18900 1620 18920 1660
rect 18960 1620 18980 1660
rect 19020 1620 19040 1660
rect 19080 1620 19100 1660
rect 18900 1600 19100 1620
rect 22500 1780 22700 11920
rect 26100 12080 26300 12100
rect 26100 12040 26120 12080
rect 26160 12040 26180 12080
rect 26220 12040 26240 12080
rect 26280 12040 26300 12080
rect 26100 12020 26300 12040
rect 26100 11980 26120 12020
rect 26160 11980 26180 12020
rect 26220 11980 26240 12020
rect 26280 11980 26300 12020
rect 26100 11960 26300 11980
rect 26100 11920 26120 11960
rect 26160 11920 26180 11960
rect 26220 11920 26240 11960
rect 26280 11920 26300 11960
rect 24300 11680 24500 11700
rect 24300 11640 24320 11680
rect 24360 11640 24380 11680
rect 24420 11640 24440 11680
rect 24480 11640 24500 11680
rect 24300 11620 24500 11640
rect 24300 11580 24320 11620
rect 24360 11580 24380 11620
rect 24420 11580 24440 11620
rect 24480 11580 24500 11620
rect 24300 11560 24500 11580
rect 24300 11520 24320 11560
rect 24360 11520 24380 11560
rect 24420 11520 24440 11560
rect 24480 11520 24500 11560
rect 24300 2180 24500 11520
rect 24300 2140 24320 2180
rect 24360 2140 24380 2180
rect 24420 2140 24440 2180
rect 24480 2140 24500 2180
rect 24300 2120 24500 2140
rect 24300 2080 24320 2120
rect 24360 2080 24380 2120
rect 24420 2080 24440 2120
rect 24480 2080 24500 2120
rect 24300 2060 24500 2080
rect 24300 2020 24320 2060
rect 24360 2020 24380 2060
rect 24420 2020 24440 2060
rect 24480 2020 24500 2060
rect 24300 2000 24500 2020
rect 22500 1740 22520 1780
rect 22560 1740 22580 1780
rect 22620 1740 22640 1780
rect 22680 1740 22700 1780
rect 22500 1720 22700 1740
rect 22500 1680 22520 1720
rect 22560 1680 22580 1720
rect 22620 1680 22640 1720
rect 22680 1680 22700 1720
rect 22500 1660 22700 1680
rect 22500 1620 22520 1660
rect 22560 1620 22580 1660
rect 22620 1620 22640 1660
rect 22680 1620 22700 1660
rect 22500 1600 22700 1620
rect 26100 1780 26300 11920
rect 29700 12080 29900 12100
rect 29700 12040 29720 12080
rect 29760 12040 29780 12080
rect 29820 12040 29840 12080
rect 29880 12040 29900 12080
rect 29700 12020 29900 12040
rect 29700 11980 29720 12020
rect 29760 11980 29780 12020
rect 29820 11980 29840 12020
rect 29880 11980 29900 12020
rect 29700 11960 29900 11980
rect 29700 11920 29720 11960
rect 29760 11920 29780 11960
rect 29820 11920 29840 11960
rect 29880 11920 29900 11960
rect 27900 11680 28100 11700
rect 27900 11640 27920 11680
rect 27960 11640 27980 11680
rect 28020 11640 28040 11680
rect 28080 11640 28100 11680
rect 27900 11620 28100 11640
rect 27900 11580 27920 11620
rect 27960 11580 27980 11620
rect 28020 11580 28040 11620
rect 28080 11580 28100 11620
rect 27900 11560 28100 11580
rect 27900 11520 27920 11560
rect 27960 11520 27980 11560
rect 28020 11520 28040 11560
rect 28080 11520 28100 11560
rect 27900 2180 28100 11520
rect 27900 2140 27920 2180
rect 27960 2140 27980 2180
rect 28020 2140 28040 2180
rect 28080 2140 28100 2180
rect 27900 2120 28100 2140
rect 27900 2080 27920 2120
rect 27960 2080 27980 2120
rect 28020 2080 28040 2120
rect 28080 2080 28100 2120
rect 27900 2060 28100 2080
rect 27900 2020 27920 2060
rect 27960 2020 27980 2060
rect 28020 2020 28040 2060
rect 28080 2020 28100 2060
rect 27900 2000 28100 2020
rect 26100 1740 26120 1780
rect 26160 1740 26180 1780
rect 26220 1740 26240 1780
rect 26280 1740 26300 1780
rect 26100 1720 26300 1740
rect 26100 1680 26120 1720
rect 26160 1680 26180 1720
rect 26220 1680 26240 1720
rect 26280 1680 26300 1720
rect 26100 1660 26300 1680
rect 26100 1620 26120 1660
rect 26160 1620 26180 1660
rect 26220 1620 26240 1660
rect 26280 1620 26300 1660
rect 26100 1600 26300 1620
rect 29700 1780 29900 11920
rect 31500 11680 31700 11700
rect 31500 11640 31520 11680
rect 31560 11640 31580 11680
rect 31620 11640 31640 11680
rect 31680 11640 31700 11680
rect 31500 11620 31700 11640
rect 31500 11580 31520 11620
rect 31560 11580 31580 11620
rect 31620 11580 31640 11620
rect 31680 11580 31700 11620
rect 31500 11560 31700 11580
rect 31500 11520 31520 11560
rect 31560 11520 31580 11560
rect 31620 11520 31640 11560
rect 31680 11520 31700 11560
rect 31500 2180 31700 11520
rect 31500 2140 31520 2180
rect 31560 2140 31580 2180
rect 31620 2140 31640 2180
rect 31680 2140 31700 2180
rect 31500 2120 31700 2140
rect 31500 2080 31520 2120
rect 31560 2080 31580 2120
rect 31620 2080 31640 2120
rect 31680 2080 31700 2120
rect 31500 2060 31700 2080
rect 31500 2020 31520 2060
rect 31560 2020 31580 2060
rect 31620 2020 31640 2060
rect 31680 2020 31700 2060
rect 31500 2000 31700 2020
rect 29700 1740 29720 1780
rect 29760 1740 29780 1780
rect 29820 1740 29840 1780
rect 29880 1740 29900 1780
rect 29700 1720 29900 1740
rect 29700 1680 29720 1720
rect 29760 1680 29780 1720
rect 29820 1680 29840 1720
rect 29880 1680 29900 1720
rect 29700 1660 29900 1680
rect 29700 1620 29720 1660
rect 29760 1620 29780 1660
rect 29820 1620 29840 1660
rect 29880 1620 29900 1660
rect 29700 1600 29900 1620
<< end >>
