magic
tech sky130A
timestamp 1637233519
<< psubdiff >>
rect 720 3630 760 3660
rect 790 3630 820 3660
rect 850 3630 880 3660
rect 910 3630 940 3660
rect 970 3630 1000 3660
rect 1030 3630 1060 3660
rect 1090 3630 1120 3660
rect 1150 3630 1180 3660
rect 1210 3630 1240 3660
rect 1270 3630 1300 3660
rect 1330 3630 1360 3660
rect 1390 3630 1420 3660
rect 1450 3630 1480 3660
rect 1510 3630 1540 3660
rect 1570 3630 1600 3660
rect 1630 3630 1660 3660
rect 1690 3630 1720 3660
rect 1750 3630 1780 3660
rect 1810 3630 1840 3660
rect 1870 3630 1900 3660
rect 1930 3630 1960 3660
rect 1990 3630 2020 3660
rect 2050 3630 2080 3660
rect 2110 3630 2140 3660
rect 2170 3630 2200 3660
rect 2230 3630 2260 3660
rect 2290 3630 2320 3660
rect 2350 3630 2380 3660
rect 2410 3630 2440 3660
rect 2470 3630 2500 3660
rect 2530 3630 2560 3660
rect 2590 3630 2620 3660
rect 2650 3630 2680 3660
rect 2710 3630 2740 3660
rect 2770 3630 2800 3660
rect 2830 3630 2860 3660
rect 2890 3630 2920 3660
rect 2950 3630 2980 3660
rect 3010 3630 3040 3660
rect 3070 3630 3100 3660
rect 3130 3630 3160 3660
rect 3190 3630 3220 3660
rect 3250 3630 3280 3660
rect 3310 3630 3340 3660
rect 3370 3630 3400 3660
rect 3430 3630 3460 3660
rect 3490 3630 3520 3660
rect 3550 3630 3580 3660
rect 3610 3630 3640 3660
rect 3670 3630 3700 3660
rect 3730 3630 3760 3660
rect 3790 3630 3820 3660
rect 3850 3630 3880 3660
rect 3910 3630 3940 3660
rect 3970 3630 4000 3660
rect 4030 3630 4060 3660
rect 4090 3630 4120 3660
rect 4150 3630 4180 3660
rect 4210 3630 4240 3660
rect 4270 3630 4300 3660
rect 4330 3630 4360 3660
rect 4390 3630 4420 3660
rect 4450 3630 4480 3660
rect 4510 3630 4540 3660
rect 4570 3630 4600 3660
rect 4630 3630 4660 3660
rect 4690 3630 4720 3660
rect 4750 3630 4780 3660
rect 4810 3630 4840 3660
rect 4870 3630 4900 3660
rect 4930 3630 4960 3660
rect 4990 3630 5020 3660
rect 5050 3630 5080 3660
rect 5110 3630 5140 3660
rect 5170 3630 5200 3660
rect 5230 3630 5260 3660
rect 5290 3630 5320 3660
rect 5350 3630 5380 3660
rect 5410 3630 5440 3660
rect 5470 3630 5500 3660
rect 5530 3630 5560 3660
rect 5590 3630 5620 3660
rect 5650 3630 5680 3660
rect 5710 3630 5740 3660
rect 5770 3630 5800 3660
rect 5830 3630 5860 3660
rect 5890 3630 5920 3660
rect 5950 3630 5980 3660
rect 6010 3630 6040 3660
rect 6070 3630 6100 3660
rect 6130 3630 6160 3660
rect 6190 3630 6220 3660
rect 6250 3630 6280 3660
rect 6310 3630 6340 3660
rect 6370 3630 6400 3660
rect 6430 3630 6460 3660
rect 6490 3630 6520 3660
rect 6550 3630 6580 3660
rect 6610 3630 6640 3660
rect 6670 3630 6700 3660
rect 6730 3630 6760 3660
rect 6790 3630 6820 3660
rect 6850 3630 6880 3660
rect 6910 3630 6940 3660
rect 6970 3630 7000 3660
rect 7030 3630 7060 3660
rect 7090 3630 7120 3660
rect 7150 3630 7180 3660
rect 7210 3630 7240 3660
rect 7270 3630 7300 3660
rect 7330 3630 7360 3660
rect 7390 3630 7420 3660
rect 7450 3630 7480 3660
rect 7510 3630 7540 3660
rect 7570 3630 7600 3660
rect 7630 3630 7660 3660
rect 7690 3630 7720 3660
rect 7750 3630 7780 3660
rect 7810 3630 7840 3660
rect 7870 3630 7900 3660
rect 7930 3630 7960 3660
rect 7990 3630 8020 3660
rect 8050 3630 8080 3660
rect 8110 3630 8140 3660
rect 8170 3630 8200 3660
rect 8230 3630 8260 3660
rect 8290 3630 8320 3660
rect 8350 3630 8380 3660
rect 8410 3630 8440 3660
rect 8470 3630 8500 3660
rect 8530 3630 8560 3660
rect 8590 3630 8620 3660
rect 8650 3630 8680 3660
rect 8710 3630 8740 3660
rect 8770 3630 8800 3660
rect 8830 3630 8860 3660
rect 8890 3630 8920 3660
rect 8950 3630 8980 3660
rect 9010 3630 9040 3660
rect 9070 3630 9100 3660
rect 9130 3630 9160 3660
rect 9190 3630 9220 3660
rect 9250 3630 9280 3660
rect 9310 3630 9340 3660
rect 9370 3630 9400 3660
rect 9430 3630 9460 3660
rect 9490 3630 9520 3660
rect 720 3610 750 3630
rect 720 3550 750 3580
rect 720 3490 750 3520
rect 720 3430 750 3460
rect 720 3370 750 3400
rect 720 3310 750 3340
rect 720 3250 750 3280
rect 720 3190 750 3220
rect 720 3130 750 3160
rect 720 3070 750 3100
rect 720 3010 750 3040
rect 720 2950 750 2980
rect 720 2890 750 2920
rect 720 2830 750 2860
rect 720 2770 750 2800
rect 720 2710 750 2740
rect 720 2650 750 2680
rect 720 2590 750 2620
rect 720 2530 750 2560
rect 720 2470 750 2500
rect 720 2410 750 2440
rect 720 2350 750 2380
rect 720 2290 750 2320
rect 720 2230 750 2260
rect 720 2170 750 2200
rect 720 2120 750 2140
rect 720 2060 750 2080
rect 720 2000 750 2020
rect 720 1940 750 1960
rect 720 1845 750 1910
rect 9550 3610 9580 3660
rect 9550 3550 9580 3580
rect 9550 3490 9580 3520
rect 9550 3430 9580 3460
rect 9550 3370 9580 3400
rect 9550 3310 9580 3340
rect 9550 3250 9580 3280
rect 9550 3190 9580 3220
rect 9550 3130 9580 3160
rect 9550 3070 9580 3100
rect 9550 3010 9580 3040
rect 9550 2950 9580 2980
rect 9550 2890 9580 2920
rect 9550 2830 9580 2860
rect 9550 2770 9580 2800
rect 9550 2710 9580 2740
rect 9550 2650 9580 2680
rect 9550 2590 9580 2620
rect 9550 2530 9580 2560
rect 9550 2470 9580 2500
rect 9550 2410 9580 2440
rect 9550 2350 9580 2380
rect 9550 2290 9580 2320
rect 9550 2230 9580 2260
rect 9550 2170 9580 2200
rect 9550 2120 9580 2140
rect 9550 2060 9580 2080
rect 9550 2000 9580 2020
rect 9550 1940 9580 1960
rect 9550 1845 9580 1910
rect 170 1787 200 1845
rect 230 1815 260 1845
rect 290 1815 320 1845
rect 350 1815 380 1845
rect 410 1815 440 1845
rect 470 1815 500 1845
rect 530 1815 560 1845
rect 590 1815 620 1845
rect 650 1815 680 1845
rect 710 1815 740 1845
rect 770 1815 800 1845
rect 830 1815 860 1845
rect 890 1815 910 1845
rect 940 1815 970 1845
rect 1000 1815 1030 1845
rect 1060 1815 1090 1845
rect 1120 1815 1150 1845
rect 1180 1815 1210 1845
rect 1240 1815 1270 1845
rect 1300 1815 1330 1845
rect 1360 1815 1390 1845
rect 1420 1815 1450 1845
rect 1480 1815 1510 1845
rect 1540 1815 1570 1845
rect 1600 1815 1630 1845
rect 1660 1815 1690 1845
rect 1720 1815 1750 1845
rect 1780 1815 1810 1845
rect 1840 1815 1870 1845
rect 1900 1815 1930 1845
rect 1960 1815 1990 1845
rect 2020 1815 2050 1845
rect 2080 1815 2110 1845
rect 2140 1815 2170 1845
rect 2200 1815 2230 1845
rect 2260 1815 2290 1845
rect 2320 1815 2350 1845
rect 2380 1815 2410 1845
rect 2440 1815 2470 1845
rect 2500 1815 2530 1845
rect 2560 1815 2590 1845
rect 2620 1815 2650 1845
rect 2680 1815 2710 1845
rect 2740 1815 2770 1845
rect 2800 1815 2830 1845
rect 2860 1815 2890 1845
rect 2920 1815 2950 1845
rect 2980 1815 3010 1845
rect 3040 1815 3070 1845
rect 3100 1815 3130 1845
rect 3160 1815 3190 1845
rect 3220 1815 3250 1845
rect 3280 1815 3310 1845
rect 3340 1815 3370 1845
rect 3400 1815 3430 1845
rect 3460 1815 3490 1845
rect 3520 1815 3550 1845
rect 3580 1815 3610 1845
rect 3640 1815 3670 1845
rect 3700 1815 3730 1845
rect 3760 1815 3790 1845
rect 3820 1815 3850 1845
rect 3880 1815 3910 1845
rect 3940 1815 3970 1845
rect 4000 1815 4030 1845
rect 4060 1815 4090 1845
rect 4120 1815 4150 1845
rect 4180 1815 4210 1845
rect 4240 1815 4270 1845
rect 4300 1815 4330 1845
rect 4360 1815 4390 1845
rect 4420 1815 4450 1845
rect 4480 1815 4510 1845
rect 4540 1815 4570 1845
rect 4600 1815 4630 1845
rect 4660 1815 4690 1845
rect 4720 1815 4750 1845
rect 4780 1815 4810 1845
rect 4840 1815 4870 1845
rect 4900 1815 4930 1845
rect 4960 1815 4990 1845
rect 5020 1815 5050 1845
rect 5080 1815 5110 1845
rect 5140 1815 5170 1845
rect 5200 1815 5230 1845
rect 5260 1815 5290 1845
rect 5320 1815 5350 1845
rect 5380 1815 5410 1845
rect 5440 1815 5470 1845
rect 5500 1815 5530 1845
rect 5560 1815 5590 1845
rect 5620 1815 5650 1845
rect 5680 1815 5710 1845
rect 5740 1815 5770 1845
rect 5800 1815 5830 1845
rect 5860 1815 5890 1845
rect 5920 1815 5950 1845
rect 5980 1815 6010 1845
rect 6040 1815 6070 1845
rect 6100 1815 6130 1845
rect 6160 1815 6190 1845
rect 6220 1815 6250 1845
rect 6280 1815 6310 1845
rect 6340 1815 6370 1845
rect 6400 1815 6430 1845
rect 6460 1815 6490 1845
rect 6520 1815 6550 1845
rect 6580 1815 6610 1845
rect 6640 1815 6670 1845
rect 6700 1815 6730 1845
rect 6760 1815 6790 1845
rect 6820 1815 6850 1845
rect 6880 1815 6910 1845
rect 6940 1815 6970 1845
rect 7000 1815 7030 1845
rect 7060 1815 7090 1845
rect 7120 1815 7150 1845
rect 7180 1815 7210 1845
rect 7240 1815 7270 1845
rect 7300 1815 7330 1845
rect 7360 1815 7390 1845
rect 7420 1815 7450 1845
rect 7480 1815 7510 1845
rect 7540 1815 7570 1845
rect 7600 1815 7630 1845
rect 7660 1815 7690 1845
rect 7720 1815 7750 1845
rect 7780 1815 7810 1845
rect 7840 1815 7870 1845
rect 7900 1815 7930 1845
rect 7960 1815 7990 1845
rect 8020 1815 8050 1845
rect 8080 1815 8110 1845
rect 8140 1815 8170 1845
rect 8200 1815 8230 1845
rect 8260 1815 8290 1845
rect 8320 1815 8350 1845
rect 8380 1815 8410 1845
rect 8440 1815 8470 1845
rect 8500 1815 8530 1845
rect 8560 1815 8590 1845
rect 8620 1815 8650 1845
rect 8680 1815 8710 1845
rect 8740 1815 8770 1845
rect 8800 1815 8830 1845
rect 8860 1815 8890 1845
rect 8920 1815 8950 1845
rect 8980 1815 9010 1845
rect 9040 1815 9070 1845
rect 9100 1815 9130 1845
rect 9160 1815 9190 1845
rect 9220 1815 9250 1845
rect 9280 1815 9310 1845
rect 9340 1815 9370 1845
rect 9400 1815 9430 1845
rect 9460 1815 9490 1845
rect 9520 1815 9550 1845
rect 9580 1815 9610 1845
rect 9640 1815 9670 1845
rect 9700 1815 9730 1845
rect 9760 1815 9790 1845
rect 9820 1815 9850 1845
rect 9880 1815 9910 1845
rect 9940 1815 9970 1845
rect 10000 1815 10030 1845
rect 10060 1815 10090 1845
rect 10120 1815 10150 1845
rect 10180 1815 10210 1845
rect 10240 1815 10270 1845
rect 10300 1815 10330 1845
rect 10360 1815 10390 1845
rect 10420 1815 10450 1845
rect 10480 1815 10510 1845
rect 10540 1815 10570 1845
rect 10600 1815 10630 1845
rect 10660 1815 10688 1845
rect 10718 1815 10730 1845
rect 170 1727 200 1757
rect 170 1667 200 1697
rect 170 1607 200 1637
rect 170 1547 200 1577
rect 170 1487 200 1517
rect 170 1427 200 1457
rect 170 1367 200 1397
rect 170 1307 200 1337
rect 170 1247 200 1277
rect 170 1187 200 1217
rect 170 1127 200 1157
rect 170 1067 200 1097
rect 170 1007 200 1037
rect 170 947 200 977
rect 170 887 200 917
rect 170 827 200 857
rect 170 767 200 797
rect 170 707 200 737
rect 170 647 200 677
rect 170 587 200 617
rect 170 527 200 557
rect 170 467 200 497
rect 170 407 200 437
rect 170 347 200 377
rect 170 290 200 317
rect 170 230 200 260
rect 170 170 200 200
rect 170 113 200 140
rect 170 30 200 83
rect 10700 1787 10730 1815
rect 10700 1727 10730 1757
rect 10700 1667 10730 1697
rect 10700 1607 10730 1637
rect 10700 1547 10730 1577
rect 10700 1487 10730 1517
rect 10700 1427 10730 1457
rect 10700 1367 10730 1397
rect 10700 1307 10730 1337
rect 10700 1247 10730 1277
rect 10700 1187 10730 1217
rect 10700 1127 10730 1157
rect 10700 1067 10730 1097
rect 10700 1007 10730 1037
rect 10700 947 10730 977
rect 10700 887 10730 917
rect 10700 827 10730 857
rect 10700 767 10730 797
rect 10700 707 10730 737
rect 10700 647 10730 677
rect 10700 587 10730 617
rect 10700 527 10730 557
rect 10700 467 10730 497
rect 10700 407 10730 437
rect 10700 347 10730 377
rect 10700 290 10730 317
rect 10700 230 10730 260
rect 10700 170 10730 200
rect 10700 113 10730 140
rect 10700 30 10730 83
rect 170 0 210 30
rect 240 0 270 30
rect 300 0 330 30
rect 360 0 390 30
rect 420 0 450 30
rect 480 0 510 30
rect 540 0 570 30
rect 600 0 630 30
rect 660 0 690 30
rect 720 0 750 30
rect 780 0 810 30
rect 840 0 870 30
rect 900 0 930 30
rect 960 0 990 30
rect 1020 0 1050 30
rect 1080 0 1110 30
rect 1140 0 1170 30
rect 1200 0 1230 30
rect 1260 0 1290 30
rect 1320 0 1350 30
rect 1380 0 1410 30
rect 1440 0 1470 30
rect 1500 0 1530 30
rect 1560 0 1590 30
rect 1620 0 1650 30
rect 1680 0 1710 30
rect 1740 0 1770 30
rect 1800 0 1830 30
rect 1860 0 1890 30
rect 1920 0 1950 30
rect 1980 0 2010 30
rect 2040 0 2070 30
rect 2100 0 2130 30
rect 2160 0 2190 30
rect 2220 0 2250 30
rect 2280 0 2310 30
rect 2340 0 2370 30
rect 2400 0 2430 30
rect 2460 0 2490 30
rect 2520 0 2550 30
rect 2580 0 2610 30
rect 2640 0 2670 30
rect 2700 0 2730 30
rect 2760 0 2790 30
rect 2820 0 2850 30
rect 2880 0 2910 30
rect 2940 0 2970 30
rect 3000 0 3030 30
rect 3060 0 3090 30
rect 3120 0 3150 30
rect 3180 0 3210 30
rect 3240 0 3270 30
rect 3300 0 3330 30
rect 3360 0 3390 30
rect 3420 0 3450 30
rect 3480 0 3510 30
rect 3540 0 3570 30
rect 3600 0 3630 30
rect 3660 0 3690 30
rect 3720 0 3750 30
rect 3780 0 3810 30
rect 3840 0 3870 30
rect 3900 0 3930 30
rect 3960 0 3990 30
rect 4020 0 4050 30
rect 4080 0 4110 30
rect 4140 0 4170 30
rect 4200 0 4230 30
rect 4260 0 4290 30
rect 4320 0 4350 30
rect 4380 0 4410 30
rect 4440 0 4470 30
rect 4500 0 4530 30
rect 4560 0 4590 30
rect 4620 0 4650 30
rect 4680 0 4710 30
rect 4740 0 4770 30
rect 4800 0 4830 30
rect 4860 0 4890 30
rect 4920 0 4950 30
rect 4980 0 5010 30
rect 5040 0 5070 30
rect 5100 0 5130 30
rect 5160 0 5190 30
rect 5220 0 5250 30
rect 5280 0 5310 30
rect 5340 0 5370 30
rect 5400 0 5430 30
rect 5460 0 5490 30
rect 5520 0 5550 30
rect 5580 0 5610 30
rect 5640 0 5670 30
rect 5700 0 5730 30
rect 5760 0 5790 30
rect 5820 0 5850 30
rect 5880 0 5910 30
rect 5940 0 5970 30
rect 6000 0 6030 30
rect 6060 0 6090 30
rect 6120 0 6150 30
rect 6180 0 6210 30
rect 6240 0 6270 30
rect 6300 0 6330 30
rect 6360 0 6390 30
rect 6420 0 6450 30
rect 6480 0 6510 30
rect 6540 0 6570 30
rect 6600 0 6630 30
rect 6660 0 6690 30
rect 6720 0 6750 30
rect 6780 0 6810 30
rect 6840 0 6870 30
rect 6900 0 6930 30
rect 6960 0 6990 30
rect 7020 0 7050 30
rect 7080 0 7110 30
rect 7140 0 7170 30
rect 7200 0 7230 30
rect 7260 0 7290 30
rect 7320 0 7350 30
rect 7380 0 7410 30
rect 7440 0 7470 30
rect 7500 0 7530 30
rect 7560 0 7590 30
rect 7620 0 7650 30
rect 7680 0 7710 30
rect 7740 0 7770 30
rect 7800 0 7830 30
rect 7860 0 7890 30
rect 7920 0 7950 30
rect 7980 0 8010 30
rect 8040 0 8070 30
rect 8100 0 8130 30
rect 8160 0 8190 30
rect 8220 0 8250 30
rect 8280 0 8310 30
rect 8340 0 8370 30
rect 8400 0 8430 30
rect 8460 0 8490 30
rect 8520 0 8550 30
rect 8580 0 8610 30
rect 8640 0 8670 30
rect 8700 0 8730 30
rect 8760 0 8790 30
rect 8820 0 8850 30
rect 8880 0 8910 30
rect 8940 0 8970 30
rect 9000 0 9030 30
rect 9060 0 9090 30
rect 9120 0 9150 30
rect 9180 0 9210 30
rect 9240 0 9270 30
rect 9300 0 9330 30
rect 9360 0 9390 30
rect 9420 0 9450 30
rect 9480 0 9510 30
rect 9540 0 9570 30
rect 9600 0 9630 30
rect 9660 0 9690 30
rect 9720 0 9750 30
rect 9780 0 9810 30
rect 9840 0 9870 30
rect 9900 0 9930 30
rect 9960 0 9990 30
rect 10020 0 10050 30
rect 10080 0 10110 30
rect 10140 0 10170 30
rect 10200 0 10230 30
rect 10260 0 10290 30
rect 10320 0 10350 30
rect 10380 0 10410 30
rect 10440 0 10470 30
rect 10500 0 10530 30
rect 10560 0 10590 30
rect 10620 0 10650 30
rect 10680 0 10730 30
<< psubdiffcont >>
rect 760 3630 790 3660
rect 820 3630 850 3660
rect 880 3630 910 3660
rect 940 3630 970 3660
rect 1000 3630 1030 3660
rect 1060 3630 1090 3660
rect 1120 3630 1150 3660
rect 1180 3630 1210 3660
rect 1240 3630 1270 3660
rect 1300 3630 1330 3660
rect 1360 3630 1390 3660
rect 1420 3630 1450 3660
rect 1480 3630 1510 3660
rect 1540 3630 1570 3660
rect 1600 3630 1630 3660
rect 1660 3630 1690 3660
rect 1720 3630 1750 3660
rect 1780 3630 1810 3660
rect 1840 3630 1870 3660
rect 1900 3630 1930 3660
rect 1960 3630 1990 3660
rect 2020 3630 2050 3660
rect 2080 3630 2110 3660
rect 2140 3630 2170 3660
rect 2200 3630 2230 3660
rect 2260 3630 2290 3660
rect 2320 3630 2350 3660
rect 2380 3630 2410 3660
rect 2440 3630 2470 3660
rect 2500 3630 2530 3660
rect 2560 3630 2590 3660
rect 2620 3630 2650 3660
rect 2680 3630 2710 3660
rect 2740 3630 2770 3660
rect 2800 3630 2830 3660
rect 2860 3630 2890 3660
rect 2920 3630 2950 3660
rect 2980 3630 3010 3660
rect 3040 3630 3070 3660
rect 3100 3630 3130 3660
rect 3160 3630 3190 3660
rect 3220 3630 3250 3660
rect 3280 3630 3310 3660
rect 3340 3630 3370 3660
rect 3400 3630 3430 3660
rect 3460 3630 3490 3660
rect 3520 3630 3550 3660
rect 3580 3630 3610 3660
rect 3640 3630 3670 3660
rect 3700 3630 3730 3660
rect 3760 3630 3790 3660
rect 3820 3630 3850 3660
rect 3880 3630 3910 3660
rect 3940 3630 3970 3660
rect 4000 3630 4030 3660
rect 4060 3630 4090 3660
rect 4120 3630 4150 3660
rect 4180 3630 4210 3660
rect 4240 3630 4270 3660
rect 4300 3630 4330 3660
rect 4360 3630 4390 3660
rect 4420 3630 4450 3660
rect 4480 3630 4510 3660
rect 4540 3630 4570 3660
rect 4600 3630 4630 3660
rect 4660 3630 4690 3660
rect 4720 3630 4750 3660
rect 4780 3630 4810 3660
rect 4840 3630 4870 3660
rect 4900 3630 4930 3660
rect 4960 3630 4990 3660
rect 5020 3630 5050 3660
rect 5080 3630 5110 3660
rect 5140 3630 5170 3660
rect 5200 3630 5230 3660
rect 5260 3630 5290 3660
rect 5320 3630 5350 3660
rect 5380 3630 5410 3660
rect 5440 3630 5470 3660
rect 5500 3630 5530 3660
rect 5560 3630 5590 3660
rect 5620 3630 5650 3660
rect 5680 3630 5710 3660
rect 5740 3630 5770 3660
rect 5800 3630 5830 3660
rect 5860 3630 5890 3660
rect 5920 3630 5950 3660
rect 5980 3630 6010 3660
rect 6040 3630 6070 3660
rect 6100 3630 6130 3660
rect 6160 3630 6190 3660
rect 6220 3630 6250 3660
rect 6280 3630 6310 3660
rect 6340 3630 6370 3660
rect 6400 3630 6430 3660
rect 6460 3630 6490 3660
rect 6520 3630 6550 3660
rect 6580 3630 6610 3660
rect 6640 3630 6670 3660
rect 6700 3630 6730 3660
rect 6760 3630 6790 3660
rect 6820 3630 6850 3660
rect 6880 3630 6910 3660
rect 6940 3630 6970 3660
rect 7000 3630 7030 3660
rect 7060 3630 7090 3660
rect 7120 3630 7150 3660
rect 7180 3630 7210 3660
rect 7240 3630 7270 3660
rect 7300 3630 7330 3660
rect 7360 3630 7390 3660
rect 7420 3630 7450 3660
rect 7480 3630 7510 3660
rect 7540 3630 7570 3660
rect 7600 3630 7630 3660
rect 7660 3630 7690 3660
rect 7720 3630 7750 3660
rect 7780 3630 7810 3660
rect 7840 3630 7870 3660
rect 7900 3630 7930 3660
rect 7960 3630 7990 3660
rect 8020 3630 8050 3660
rect 8080 3630 8110 3660
rect 8140 3630 8170 3660
rect 8200 3630 8230 3660
rect 8260 3630 8290 3660
rect 8320 3630 8350 3660
rect 8380 3630 8410 3660
rect 8440 3630 8470 3660
rect 8500 3630 8530 3660
rect 8560 3630 8590 3660
rect 8620 3630 8650 3660
rect 8680 3630 8710 3660
rect 8740 3630 8770 3660
rect 8800 3630 8830 3660
rect 8860 3630 8890 3660
rect 8920 3630 8950 3660
rect 8980 3630 9010 3660
rect 9040 3630 9070 3660
rect 9100 3630 9130 3660
rect 9160 3630 9190 3660
rect 9220 3630 9250 3660
rect 9280 3630 9310 3660
rect 9340 3630 9370 3660
rect 9400 3630 9430 3660
rect 9460 3630 9490 3660
rect 9520 3630 9550 3660
rect 720 3580 750 3610
rect 720 3520 750 3550
rect 720 3460 750 3490
rect 720 3400 750 3430
rect 720 3340 750 3370
rect 720 3280 750 3310
rect 720 3220 750 3250
rect 720 3160 750 3190
rect 720 3100 750 3130
rect 720 3040 750 3070
rect 720 2980 750 3010
rect 720 2920 750 2950
rect 720 2860 750 2890
rect 720 2800 750 2830
rect 720 2740 750 2770
rect 720 2680 750 2710
rect 720 2620 750 2650
rect 720 2560 750 2590
rect 720 2500 750 2530
rect 720 2440 750 2470
rect 720 2380 750 2410
rect 720 2320 750 2350
rect 720 2260 750 2290
rect 720 2200 750 2230
rect 720 2140 750 2170
rect 720 2080 750 2120
rect 720 2020 750 2060
rect 720 1960 750 2000
rect 720 1910 750 1940
rect 9550 3580 9580 3610
rect 9550 3520 9580 3550
rect 9550 3460 9580 3490
rect 9550 3400 9580 3430
rect 9550 3340 9580 3370
rect 9550 3280 9580 3310
rect 9550 3220 9580 3250
rect 9550 3160 9580 3190
rect 9550 3100 9580 3130
rect 9550 3040 9580 3070
rect 9550 2980 9580 3010
rect 9550 2920 9580 2950
rect 9550 2860 9580 2890
rect 9550 2800 9580 2830
rect 9550 2740 9580 2770
rect 9550 2680 9580 2710
rect 9550 2620 9580 2650
rect 9550 2560 9580 2590
rect 9550 2500 9580 2530
rect 9550 2440 9580 2470
rect 9550 2380 9580 2410
rect 9550 2320 9580 2350
rect 9550 2260 9580 2290
rect 9550 2200 9580 2230
rect 9550 2140 9580 2170
rect 9550 2080 9580 2120
rect 9550 2020 9580 2060
rect 9550 1960 9580 2000
rect 9550 1910 9580 1940
rect 200 1815 230 1845
rect 260 1815 290 1845
rect 320 1815 350 1845
rect 380 1815 410 1845
rect 440 1815 470 1845
rect 500 1815 530 1845
rect 560 1815 590 1845
rect 620 1815 650 1845
rect 680 1815 710 1845
rect 740 1815 770 1845
rect 800 1815 830 1845
rect 860 1815 890 1845
rect 910 1815 940 1845
rect 970 1815 1000 1845
rect 1030 1815 1060 1845
rect 1090 1815 1120 1845
rect 1150 1815 1180 1845
rect 1210 1815 1240 1845
rect 1270 1815 1300 1845
rect 1330 1815 1360 1845
rect 1390 1815 1420 1845
rect 1450 1815 1480 1845
rect 1510 1815 1540 1845
rect 1570 1815 1600 1845
rect 1630 1815 1660 1845
rect 1690 1815 1720 1845
rect 1750 1815 1780 1845
rect 1810 1815 1840 1845
rect 1870 1815 1900 1845
rect 1930 1815 1960 1845
rect 1990 1815 2020 1845
rect 2050 1815 2080 1845
rect 2110 1815 2140 1845
rect 2170 1815 2200 1845
rect 2230 1815 2260 1845
rect 2290 1815 2320 1845
rect 2350 1815 2380 1845
rect 2410 1815 2440 1845
rect 2470 1815 2500 1845
rect 2530 1815 2560 1845
rect 2590 1815 2620 1845
rect 2650 1815 2680 1845
rect 2710 1815 2740 1845
rect 2770 1815 2800 1845
rect 2830 1815 2860 1845
rect 2890 1815 2920 1845
rect 2950 1815 2980 1845
rect 3010 1815 3040 1845
rect 3070 1815 3100 1845
rect 3130 1815 3160 1845
rect 3190 1815 3220 1845
rect 3250 1815 3280 1845
rect 3310 1815 3340 1845
rect 3370 1815 3400 1845
rect 3430 1815 3460 1845
rect 3490 1815 3520 1845
rect 3550 1815 3580 1845
rect 3610 1815 3640 1845
rect 3670 1815 3700 1845
rect 3730 1815 3760 1845
rect 3790 1815 3820 1845
rect 3850 1815 3880 1845
rect 3910 1815 3940 1845
rect 3970 1815 4000 1845
rect 4030 1815 4060 1845
rect 4090 1815 4120 1845
rect 4150 1815 4180 1845
rect 4210 1815 4240 1845
rect 4270 1815 4300 1845
rect 4330 1815 4360 1845
rect 4390 1815 4420 1845
rect 4450 1815 4480 1845
rect 4510 1815 4540 1845
rect 4570 1815 4600 1845
rect 4630 1815 4660 1845
rect 4690 1815 4720 1845
rect 4750 1815 4780 1845
rect 4810 1815 4840 1845
rect 4870 1815 4900 1845
rect 4930 1815 4960 1845
rect 4990 1815 5020 1845
rect 5050 1815 5080 1845
rect 5110 1815 5140 1845
rect 5170 1815 5200 1845
rect 5230 1815 5260 1845
rect 5290 1815 5320 1845
rect 5350 1815 5380 1845
rect 5410 1815 5440 1845
rect 5470 1815 5500 1845
rect 5530 1815 5560 1845
rect 5590 1815 5620 1845
rect 5650 1815 5680 1845
rect 5710 1815 5740 1845
rect 5770 1815 5800 1845
rect 5830 1815 5860 1845
rect 5890 1815 5920 1845
rect 5950 1815 5980 1845
rect 6010 1815 6040 1845
rect 6070 1815 6100 1845
rect 6130 1815 6160 1845
rect 6190 1815 6220 1845
rect 6250 1815 6280 1845
rect 6310 1815 6340 1845
rect 6370 1815 6400 1845
rect 6430 1815 6460 1845
rect 6490 1815 6520 1845
rect 6550 1815 6580 1845
rect 6610 1815 6640 1845
rect 6670 1815 6700 1845
rect 6730 1815 6760 1845
rect 6790 1815 6820 1845
rect 6850 1815 6880 1845
rect 6910 1815 6940 1845
rect 6970 1815 7000 1845
rect 7030 1815 7060 1845
rect 7090 1815 7120 1845
rect 7150 1815 7180 1845
rect 7210 1815 7240 1845
rect 7270 1815 7300 1845
rect 7330 1815 7360 1845
rect 7390 1815 7420 1845
rect 7450 1815 7480 1845
rect 7510 1815 7540 1845
rect 7570 1815 7600 1845
rect 7630 1815 7660 1845
rect 7690 1815 7720 1845
rect 7750 1815 7780 1845
rect 7810 1815 7840 1845
rect 7870 1815 7900 1845
rect 7930 1815 7960 1845
rect 7990 1815 8020 1845
rect 8050 1815 8080 1845
rect 8110 1815 8140 1845
rect 8170 1815 8200 1845
rect 8230 1815 8260 1845
rect 8290 1815 8320 1845
rect 8350 1815 8380 1845
rect 8410 1815 8440 1845
rect 8470 1815 8500 1845
rect 8530 1815 8560 1845
rect 8590 1815 8620 1845
rect 8650 1815 8680 1845
rect 8710 1815 8740 1845
rect 8770 1815 8800 1845
rect 8830 1815 8860 1845
rect 8890 1815 8920 1845
rect 8950 1815 8980 1845
rect 9010 1815 9040 1845
rect 9070 1815 9100 1845
rect 9130 1815 9160 1845
rect 9190 1815 9220 1845
rect 9250 1815 9280 1845
rect 9310 1815 9340 1845
rect 9370 1815 9400 1845
rect 9430 1815 9460 1845
rect 9490 1815 9520 1845
rect 9550 1815 9580 1845
rect 9610 1815 9640 1845
rect 9670 1815 9700 1845
rect 9730 1815 9760 1845
rect 9790 1815 9820 1845
rect 9850 1815 9880 1845
rect 9910 1815 9940 1845
rect 9970 1815 10000 1845
rect 10030 1815 10060 1845
rect 10090 1815 10120 1845
rect 10150 1815 10180 1845
rect 10210 1815 10240 1845
rect 10270 1815 10300 1845
rect 10330 1815 10360 1845
rect 10390 1815 10420 1845
rect 10450 1815 10480 1845
rect 10510 1815 10540 1845
rect 10570 1815 10600 1845
rect 10630 1815 10660 1845
rect 10688 1815 10718 1845
rect 170 1757 200 1787
rect 170 1697 200 1727
rect 170 1637 200 1667
rect 170 1577 200 1607
rect 170 1517 200 1547
rect 170 1457 200 1487
rect 170 1397 200 1427
rect 170 1337 200 1367
rect 170 1277 200 1307
rect 170 1217 200 1247
rect 170 1157 200 1187
rect 170 1097 200 1127
rect 170 1037 200 1067
rect 170 977 200 1007
rect 170 917 200 947
rect 170 857 200 887
rect 170 797 200 827
rect 170 737 200 767
rect 170 677 200 707
rect 170 617 200 647
rect 170 557 200 587
rect 170 497 200 527
rect 170 437 200 467
rect 170 377 200 407
rect 170 317 200 347
rect 170 260 200 290
rect 170 200 200 230
rect 170 140 200 170
rect 170 83 200 113
rect 10700 1757 10730 1787
rect 10700 1697 10730 1727
rect 10700 1637 10730 1667
rect 10700 1577 10730 1607
rect 10700 1517 10730 1547
rect 10700 1457 10730 1487
rect 10700 1397 10730 1427
rect 10700 1337 10730 1367
rect 10700 1277 10730 1307
rect 10700 1217 10730 1247
rect 10700 1157 10730 1187
rect 10700 1097 10730 1127
rect 10700 1037 10730 1067
rect 10700 977 10730 1007
rect 10700 917 10730 947
rect 10700 857 10730 887
rect 10700 797 10730 827
rect 10700 737 10730 767
rect 10700 677 10730 707
rect 10700 617 10730 647
rect 10700 557 10730 587
rect 10700 497 10730 527
rect 10700 437 10730 467
rect 10700 377 10730 407
rect 10700 317 10730 347
rect 10700 260 10730 290
rect 10700 200 10730 230
rect 10700 140 10730 170
rect 10700 83 10730 113
rect 210 0 240 30
rect 270 0 300 30
rect 330 0 360 30
rect 390 0 420 30
rect 450 0 480 30
rect 510 0 540 30
rect 570 0 600 30
rect 630 0 660 30
rect 690 0 720 30
rect 750 0 780 30
rect 810 0 840 30
rect 870 0 900 30
rect 930 0 960 30
rect 990 0 1020 30
rect 1050 0 1080 30
rect 1110 0 1140 30
rect 1170 0 1200 30
rect 1230 0 1260 30
rect 1290 0 1320 30
rect 1350 0 1380 30
rect 1410 0 1440 30
rect 1470 0 1500 30
rect 1530 0 1560 30
rect 1590 0 1620 30
rect 1650 0 1680 30
rect 1710 0 1740 30
rect 1770 0 1800 30
rect 1830 0 1860 30
rect 1890 0 1920 30
rect 1950 0 1980 30
rect 2010 0 2040 30
rect 2070 0 2100 30
rect 2130 0 2160 30
rect 2190 0 2220 30
rect 2250 0 2280 30
rect 2310 0 2340 30
rect 2370 0 2400 30
rect 2430 0 2460 30
rect 2490 0 2520 30
rect 2550 0 2580 30
rect 2610 0 2640 30
rect 2670 0 2700 30
rect 2730 0 2760 30
rect 2790 0 2820 30
rect 2850 0 2880 30
rect 2910 0 2940 30
rect 2970 0 3000 30
rect 3030 0 3060 30
rect 3090 0 3120 30
rect 3150 0 3180 30
rect 3210 0 3240 30
rect 3270 0 3300 30
rect 3330 0 3360 30
rect 3390 0 3420 30
rect 3450 0 3480 30
rect 3510 0 3540 30
rect 3570 0 3600 30
rect 3630 0 3660 30
rect 3690 0 3720 30
rect 3750 0 3780 30
rect 3810 0 3840 30
rect 3870 0 3900 30
rect 3930 0 3960 30
rect 3990 0 4020 30
rect 4050 0 4080 30
rect 4110 0 4140 30
rect 4170 0 4200 30
rect 4230 0 4260 30
rect 4290 0 4320 30
rect 4350 0 4380 30
rect 4410 0 4440 30
rect 4470 0 4500 30
rect 4530 0 4560 30
rect 4590 0 4620 30
rect 4650 0 4680 30
rect 4710 0 4740 30
rect 4770 0 4800 30
rect 4830 0 4860 30
rect 4890 0 4920 30
rect 4950 0 4980 30
rect 5010 0 5040 30
rect 5070 0 5100 30
rect 5130 0 5160 30
rect 5190 0 5220 30
rect 5250 0 5280 30
rect 5310 0 5340 30
rect 5370 0 5400 30
rect 5430 0 5460 30
rect 5490 0 5520 30
rect 5550 0 5580 30
rect 5610 0 5640 30
rect 5670 0 5700 30
rect 5730 0 5760 30
rect 5790 0 5820 30
rect 5850 0 5880 30
rect 5910 0 5940 30
rect 5970 0 6000 30
rect 6030 0 6060 30
rect 6090 0 6120 30
rect 6150 0 6180 30
rect 6210 0 6240 30
rect 6270 0 6300 30
rect 6330 0 6360 30
rect 6390 0 6420 30
rect 6450 0 6480 30
rect 6510 0 6540 30
rect 6570 0 6600 30
rect 6630 0 6660 30
rect 6690 0 6720 30
rect 6750 0 6780 30
rect 6810 0 6840 30
rect 6870 0 6900 30
rect 6930 0 6960 30
rect 6990 0 7020 30
rect 7050 0 7080 30
rect 7110 0 7140 30
rect 7170 0 7200 30
rect 7230 0 7260 30
rect 7290 0 7320 30
rect 7350 0 7380 30
rect 7410 0 7440 30
rect 7470 0 7500 30
rect 7530 0 7560 30
rect 7590 0 7620 30
rect 7650 0 7680 30
rect 7710 0 7740 30
rect 7770 0 7800 30
rect 7830 0 7860 30
rect 7890 0 7920 30
rect 7950 0 7980 30
rect 8010 0 8040 30
rect 8070 0 8100 30
rect 8130 0 8160 30
rect 8190 0 8220 30
rect 8250 0 8280 30
rect 8310 0 8340 30
rect 8370 0 8400 30
rect 8430 0 8460 30
rect 8490 0 8520 30
rect 8550 0 8580 30
rect 8610 0 8640 30
rect 8670 0 8700 30
rect 8730 0 8760 30
rect 8790 0 8820 30
rect 8850 0 8880 30
rect 8910 0 8940 30
rect 8970 0 9000 30
rect 9030 0 9060 30
rect 9090 0 9120 30
rect 9150 0 9180 30
rect 9210 0 9240 30
rect 9270 0 9300 30
rect 9330 0 9360 30
rect 9390 0 9420 30
rect 9450 0 9480 30
rect 9510 0 9540 30
rect 9570 0 9600 30
rect 9630 0 9660 30
rect 9690 0 9720 30
rect 9750 0 9780 30
rect 9810 0 9840 30
rect 9870 0 9900 30
rect 9930 0 9960 30
rect 9990 0 10020 30
rect 10050 0 10080 30
rect 10110 0 10140 30
rect 10170 0 10200 30
rect 10230 0 10260 30
rect 10290 0 10320 30
rect 10350 0 10380 30
rect 10410 0 10440 30
rect 10470 0 10500 30
rect 10530 0 10560 30
rect 10590 0 10620 30
rect 10650 0 10680 30
<< locali >>
rect 720 3630 760 3660
rect 790 3630 820 3660
rect 850 3630 880 3660
rect 910 3630 940 3660
rect 970 3630 1000 3660
rect 1030 3630 1060 3660
rect 1090 3630 1120 3660
rect 1150 3630 1180 3660
rect 1210 3630 1240 3660
rect 1270 3630 1300 3660
rect 1330 3630 1360 3660
rect 1390 3630 1420 3660
rect 1450 3630 1480 3660
rect 1510 3630 1540 3660
rect 1570 3630 1600 3660
rect 1630 3630 1660 3660
rect 1690 3630 1720 3660
rect 1750 3630 1780 3660
rect 1810 3630 1840 3660
rect 1870 3630 1900 3660
rect 1930 3630 1960 3660
rect 1990 3630 2020 3660
rect 2050 3630 2080 3660
rect 2110 3630 2140 3660
rect 2170 3630 2200 3660
rect 2230 3630 2260 3660
rect 2290 3630 2320 3660
rect 2350 3630 2380 3660
rect 2410 3630 2440 3660
rect 2470 3630 2500 3660
rect 2530 3630 2560 3660
rect 2590 3630 2620 3660
rect 2650 3630 2680 3660
rect 2710 3630 2740 3660
rect 2770 3630 2800 3660
rect 2830 3630 2860 3660
rect 2890 3630 2920 3660
rect 2950 3630 2980 3660
rect 3010 3630 3040 3660
rect 3070 3630 3100 3660
rect 3130 3630 3160 3660
rect 3190 3630 3220 3660
rect 3250 3630 3280 3660
rect 3310 3630 3340 3660
rect 3370 3630 3400 3660
rect 3430 3630 3460 3660
rect 3490 3630 3520 3660
rect 3550 3630 3580 3660
rect 3610 3630 3640 3660
rect 3670 3630 3700 3660
rect 3730 3630 3760 3660
rect 3790 3630 3820 3660
rect 3850 3630 3880 3660
rect 3910 3630 3940 3660
rect 3970 3630 4000 3660
rect 4030 3630 4060 3660
rect 4090 3630 4120 3660
rect 4150 3630 4180 3660
rect 4210 3630 4240 3660
rect 4270 3630 4300 3660
rect 4330 3630 4360 3660
rect 4390 3630 4420 3660
rect 4450 3630 4480 3660
rect 4510 3630 4540 3660
rect 4570 3630 4600 3660
rect 4630 3630 4660 3660
rect 4690 3630 4720 3660
rect 4750 3630 4780 3660
rect 4810 3630 4840 3660
rect 4870 3630 4900 3660
rect 4930 3630 4960 3660
rect 4990 3630 5020 3660
rect 5050 3630 5080 3660
rect 5110 3630 5140 3660
rect 5170 3630 5200 3660
rect 5230 3630 5260 3660
rect 5290 3630 5320 3660
rect 5350 3630 5380 3660
rect 5410 3630 5440 3660
rect 5470 3630 5500 3660
rect 5530 3630 5560 3660
rect 5590 3630 5620 3660
rect 5650 3630 5680 3660
rect 5710 3630 5740 3660
rect 5770 3630 5800 3660
rect 5830 3630 5860 3660
rect 5890 3630 5920 3660
rect 5950 3630 5980 3660
rect 6010 3630 6040 3660
rect 6070 3630 6100 3660
rect 6130 3630 6160 3660
rect 6190 3630 6220 3660
rect 6250 3630 6280 3660
rect 6310 3630 6340 3660
rect 6370 3630 6400 3660
rect 6430 3630 6460 3660
rect 6490 3630 6520 3660
rect 6550 3630 6580 3660
rect 6610 3630 6640 3660
rect 6670 3630 6700 3660
rect 6730 3630 6760 3660
rect 6790 3630 6820 3660
rect 6850 3630 6880 3660
rect 6910 3630 6940 3660
rect 6970 3630 7000 3660
rect 7030 3630 7060 3660
rect 7090 3630 7120 3660
rect 7150 3630 7180 3660
rect 7210 3630 7240 3660
rect 7270 3630 7300 3660
rect 7330 3630 7360 3660
rect 7390 3630 7420 3660
rect 7450 3630 7480 3660
rect 7510 3630 7540 3660
rect 7570 3630 7600 3660
rect 7630 3630 7660 3660
rect 7690 3630 7720 3660
rect 7750 3630 7780 3660
rect 7810 3630 7840 3660
rect 7870 3630 7900 3660
rect 7930 3630 7960 3660
rect 7990 3630 8020 3660
rect 8050 3630 8080 3660
rect 8110 3630 8140 3660
rect 8170 3630 8200 3660
rect 8230 3630 8260 3660
rect 8290 3630 8320 3660
rect 8350 3630 8380 3660
rect 8410 3630 8440 3660
rect 8470 3630 8500 3660
rect 8530 3630 8560 3660
rect 8590 3630 8620 3660
rect 8650 3630 8680 3660
rect 8710 3630 8740 3660
rect 8770 3630 8800 3660
rect 8830 3630 8860 3660
rect 8890 3630 8920 3660
rect 8950 3630 8980 3660
rect 9010 3630 9040 3660
rect 9070 3630 9100 3660
rect 9130 3630 9160 3660
rect 9190 3630 9220 3660
rect 9250 3630 9280 3660
rect 9310 3630 9340 3660
rect 9370 3630 9400 3660
rect 9430 3630 9460 3660
rect 9490 3630 9520 3660
rect 720 3610 750 3630
rect 720 3550 750 3580
rect 720 3490 750 3520
rect 720 3430 750 3460
rect 720 3370 750 3400
rect 720 3310 750 3340
rect 720 3250 750 3280
rect 720 3190 750 3220
rect 720 3130 750 3160
rect 720 3070 750 3100
rect 720 3010 750 3040
rect 720 2950 750 2980
rect 720 2890 750 2920
rect 720 2830 750 2860
rect 720 2770 750 2800
rect 720 2710 750 2740
rect 720 2650 750 2680
rect 720 2590 750 2620
rect 720 2530 750 2560
rect 720 2470 750 2500
rect 720 2410 750 2440
rect 720 2350 750 2380
rect 720 2290 750 2320
rect 720 2230 750 2260
rect 720 2170 750 2200
rect 720 2120 750 2140
rect 720 2060 750 2080
rect 720 2000 750 2020
rect 720 1940 750 1960
rect 720 1845 750 1910
rect 9550 3610 9580 3660
rect 9550 3550 9580 3580
rect 9550 3490 9580 3520
rect 9550 3430 9580 3460
rect 9550 3370 9580 3400
rect 9550 3310 9580 3340
rect 9550 3250 9580 3280
rect 9550 3190 9580 3220
rect 9550 3130 9580 3160
rect 9550 3070 9580 3100
rect 9550 3010 9580 3040
rect 9550 2950 9580 2980
rect 9550 2890 9580 2920
rect 9550 2830 9580 2860
rect 9550 2770 9580 2800
rect 9550 2710 9580 2740
rect 9550 2650 9580 2680
rect 9550 2590 9580 2620
rect 9550 2530 9580 2560
rect 9550 2470 9580 2500
rect 9550 2410 9580 2440
rect 9550 2350 9580 2380
rect 9550 2290 9580 2320
rect 9550 2230 9580 2260
rect 9550 2170 9580 2200
rect 9550 2120 9580 2140
rect 9550 2060 9580 2080
rect 9550 2000 9580 2020
rect 9550 1940 9580 1960
rect 9550 1845 9580 1910
rect 170 1787 200 1845
rect 230 1815 260 1845
rect 290 1815 320 1845
rect 350 1815 380 1845
rect 410 1815 440 1845
rect 470 1815 500 1845
rect 530 1815 560 1845
rect 590 1815 620 1845
rect 650 1815 680 1845
rect 710 1815 740 1845
rect 770 1815 800 1845
rect 830 1815 860 1845
rect 890 1815 910 1845
rect 940 1815 970 1845
rect 1000 1815 1030 1845
rect 1060 1815 1090 1845
rect 1120 1815 1150 1845
rect 1180 1815 1210 1845
rect 1240 1815 1270 1845
rect 1300 1815 1330 1845
rect 1360 1815 1390 1845
rect 1420 1815 1450 1845
rect 1480 1815 1510 1845
rect 1540 1815 1570 1845
rect 1600 1815 1630 1845
rect 1660 1815 1690 1845
rect 1720 1815 1750 1845
rect 1780 1815 1810 1845
rect 1840 1815 1870 1845
rect 1900 1815 1930 1845
rect 1960 1815 1990 1845
rect 2020 1815 2050 1845
rect 2080 1815 2110 1845
rect 2140 1815 2170 1845
rect 2200 1815 2230 1845
rect 2260 1815 2290 1845
rect 2320 1815 2350 1845
rect 2380 1815 2410 1845
rect 2440 1815 2470 1845
rect 2500 1815 2530 1845
rect 2560 1815 2590 1845
rect 2620 1815 2650 1845
rect 2680 1815 2710 1845
rect 2740 1815 2770 1845
rect 2800 1815 2830 1845
rect 2860 1815 2890 1845
rect 2920 1815 2950 1845
rect 2980 1815 3010 1845
rect 3040 1815 3070 1845
rect 3100 1815 3130 1845
rect 3160 1815 3190 1845
rect 3220 1815 3250 1845
rect 3280 1815 3310 1845
rect 3340 1815 3370 1845
rect 3400 1815 3430 1845
rect 3460 1815 3490 1845
rect 3520 1815 3550 1845
rect 3580 1815 3610 1845
rect 3640 1815 3670 1845
rect 3700 1815 3730 1845
rect 3760 1815 3790 1845
rect 3820 1815 3850 1845
rect 3880 1815 3910 1845
rect 3940 1815 3970 1845
rect 4000 1815 4030 1845
rect 4060 1815 4090 1845
rect 4120 1815 4150 1845
rect 4180 1815 4210 1845
rect 4240 1815 4270 1845
rect 4300 1815 4330 1845
rect 4360 1815 4390 1845
rect 4420 1815 4450 1845
rect 4480 1815 4510 1845
rect 4540 1815 4570 1845
rect 4600 1815 4630 1845
rect 4660 1815 4690 1845
rect 4720 1815 4750 1845
rect 4780 1815 4810 1845
rect 4840 1815 4870 1845
rect 4900 1815 4930 1845
rect 4960 1815 4990 1845
rect 5020 1815 5050 1845
rect 5080 1815 5110 1845
rect 5140 1815 5170 1845
rect 5200 1815 5230 1845
rect 5260 1815 5290 1845
rect 5320 1815 5350 1845
rect 5380 1815 5410 1845
rect 5440 1815 5470 1845
rect 5500 1815 5530 1845
rect 5560 1815 5590 1845
rect 5620 1815 5650 1845
rect 5680 1815 5710 1845
rect 5740 1815 5770 1845
rect 5800 1815 5830 1845
rect 5860 1815 5890 1845
rect 5920 1815 5950 1845
rect 5980 1815 6010 1845
rect 6040 1815 6070 1845
rect 6100 1815 6130 1845
rect 6160 1815 6190 1845
rect 6220 1815 6250 1845
rect 6280 1815 6310 1845
rect 6340 1815 6370 1845
rect 6400 1815 6430 1845
rect 6460 1815 6490 1845
rect 6520 1815 6550 1845
rect 6580 1815 6610 1845
rect 6640 1815 6670 1845
rect 6700 1815 6730 1845
rect 6760 1815 6790 1845
rect 6820 1815 6850 1845
rect 6880 1815 6910 1845
rect 6940 1815 6970 1845
rect 7000 1815 7030 1845
rect 7060 1815 7090 1845
rect 7120 1815 7150 1845
rect 7180 1815 7210 1845
rect 7240 1815 7270 1845
rect 7300 1815 7330 1845
rect 7360 1815 7390 1845
rect 7420 1815 7450 1845
rect 7480 1815 7510 1845
rect 7540 1815 7570 1845
rect 7600 1815 7630 1845
rect 7660 1815 7690 1845
rect 7720 1815 7750 1845
rect 7780 1815 7810 1845
rect 7840 1815 7870 1845
rect 7900 1815 7930 1845
rect 7960 1815 7990 1845
rect 8020 1815 8050 1845
rect 8080 1815 8110 1845
rect 8140 1815 8170 1845
rect 8200 1815 8230 1845
rect 8260 1815 8290 1845
rect 8320 1815 8350 1845
rect 8380 1815 8410 1845
rect 8440 1815 8470 1845
rect 8500 1815 8530 1845
rect 8560 1815 8590 1845
rect 8620 1815 8650 1845
rect 8680 1815 8710 1845
rect 8740 1815 8770 1845
rect 8800 1815 8830 1845
rect 8860 1815 8890 1845
rect 8920 1815 8950 1845
rect 8980 1815 9010 1845
rect 9040 1815 9070 1845
rect 9100 1815 9130 1845
rect 9160 1815 9190 1845
rect 9220 1815 9250 1845
rect 9280 1815 9310 1845
rect 9340 1815 9370 1845
rect 9400 1815 9430 1845
rect 9460 1815 9490 1845
rect 9520 1815 9550 1845
rect 9580 1815 9610 1845
rect 9640 1815 9670 1845
rect 9700 1815 9730 1845
rect 9760 1815 9790 1845
rect 9820 1815 9850 1845
rect 9880 1815 9910 1845
rect 9940 1815 9970 1845
rect 10000 1815 10030 1845
rect 10060 1815 10090 1845
rect 10120 1815 10150 1845
rect 10180 1815 10210 1845
rect 10240 1815 10270 1845
rect 10300 1815 10330 1845
rect 10360 1815 10390 1845
rect 10420 1815 10450 1845
rect 10480 1815 10510 1845
rect 10540 1815 10570 1845
rect 10600 1815 10630 1845
rect 10660 1815 10688 1845
rect 10718 1815 10730 1845
rect 170 1727 200 1757
rect 170 1667 200 1697
rect 170 1607 200 1637
rect 170 1547 200 1577
rect 170 1487 200 1517
rect 170 1427 200 1457
rect 170 1367 200 1397
rect 170 1307 200 1337
rect 170 1247 200 1277
rect 170 1187 200 1217
rect 170 1127 200 1157
rect 170 1067 200 1097
rect 170 1007 200 1037
rect 170 947 200 977
rect 170 887 200 917
rect 170 827 200 857
rect 170 767 200 797
rect 170 707 200 737
rect 170 647 200 677
rect 170 587 200 617
rect 170 527 200 557
rect 170 467 200 497
rect 170 407 200 437
rect 170 347 200 377
rect 170 290 200 317
rect 170 230 200 260
rect 170 170 200 200
rect 170 113 200 140
rect 170 30 200 83
rect 10700 1787 10730 1815
rect 10700 1727 10730 1757
rect 10700 1667 10730 1697
rect 10700 1607 10730 1637
rect 10700 1547 10730 1577
rect 10700 1487 10730 1517
rect 10700 1427 10730 1457
rect 10700 1367 10730 1397
rect 10700 1307 10730 1337
rect 10700 1247 10730 1277
rect 10700 1187 10730 1217
rect 10700 1127 10730 1157
rect 10700 1067 10730 1097
rect 10700 1007 10730 1037
rect 10700 947 10730 977
rect 10700 887 10730 917
rect 10700 827 10730 857
rect 10700 767 10730 797
rect 10700 707 10730 737
rect 10700 647 10730 677
rect 10700 587 10730 617
rect 10700 527 10730 557
rect 10700 467 10730 497
rect 10700 407 10730 437
rect 10700 347 10730 377
rect 10700 290 10730 317
rect 10700 230 10730 260
rect 10700 170 10730 200
rect 10700 113 10730 140
rect 10700 30 10730 83
rect 170 0 210 30
rect 240 0 270 30
rect 300 0 330 30
rect 360 0 390 30
rect 420 0 450 30
rect 480 0 510 30
rect 540 0 570 30
rect 600 0 630 30
rect 660 0 690 30
rect 720 0 750 30
rect 780 0 810 30
rect 840 0 870 30
rect 900 0 930 30
rect 960 0 990 30
rect 1020 0 1050 30
rect 1080 0 1110 30
rect 1140 0 1170 30
rect 1200 0 1230 30
rect 1260 0 1290 30
rect 1320 0 1350 30
rect 1380 0 1410 30
rect 1440 0 1470 30
rect 1500 0 1530 30
rect 1560 0 1590 30
rect 1620 0 1650 30
rect 1680 0 1710 30
rect 1740 0 1770 30
rect 1800 0 1830 30
rect 1860 0 1890 30
rect 1920 0 1950 30
rect 1980 0 2010 30
rect 2040 0 2070 30
rect 2100 0 2130 30
rect 2160 0 2190 30
rect 2220 0 2250 30
rect 2280 0 2310 30
rect 2340 0 2370 30
rect 2400 0 2430 30
rect 2460 0 2490 30
rect 2520 0 2550 30
rect 2580 0 2610 30
rect 2640 0 2670 30
rect 2700 0 2730 30
rect 2760 0 2790 30
rect 2820 0 2850 30
rect 2880 0 2910 30
rect 2940 0 2970 30
rect 3000 0 3030 30
rect 3060 0 3090 30
rect 3120 0 3150 30
rect 3180 0 3210 30
rect 3240 0 3270 30
rect 3300 0 3330 30
rect 3360 0 3390 30
rect 3420 0 3450 30
rect 3480 0 3510 30
rect 3540 0 3570 30
rect 3600 0 3630 30
rect 3660 0 3690 30
rect 3720 0 3750 30
rect 3780 0 3810 30
rect 3840 0 3870 30
rect 3900 0 3930 30
rect 3960 0 3990 30
rect 4020 0 4050 30
rect 4080 0 4110 30
rect 4140 0 4170 30
rect 4200 0 4230 30
rect 4260 0 4290 30
rect 4320 0 4350 30
rect 4380 0 4410 30
rect 4440 0 4470 30
rect 4500 0 4530 30
rect 4560 0 4590 30
rect 4620 0 4650 30
rect 4680 0 4710 30
rect 4740 0 4770 30
rect 4800 0 4830 30
rect 4860 0 4890 30
rect 4920 0 4950 30
rect 4980 0 5010 30
rect 5040 0 5070 30
rect 5100 0 5130 30
rect 5160 0 5190 30
rect 5220 0 5250 30
rect 5280 0 5310 30
rect 5340 0 5370 30
rect 5400 0 5430 30
rect 5460 0 5490 30
rect 5520 0 5550 30
rect 5580 0 5610 30
rect 5640 0 5670 30
rect 5700 0 5730 30
rect 5760 0 5790 30
rect 5820 0 5850 30
rect 5880 0 5910 30
rect 5940 0 5970 30
rect 6000 0 6030 30
rect 6060 0 6090 30
rect 6120 0 6150 30
rect 6180 0 6210 30
rect 6240 0 6270 30
rect 6300 0 6330 30
rect 6360 0 6390 30
rect 6420 0 6450 30
rect 6480 0 6510 30
rect 6540 0 6570 30
rect 6600 0 6630 30
rect 6660 0 6690 30
rect 6720 0 6750 30
rect 6780 0 6810 30
rect 6840 0 6870 30
rect 6900 0 6930 30
rect 6960 0 6990 30
rect 7020 0 7050 30
rect 7080 0 7110 30
rect 7140 0 7170 30
rect 7200 0 7230 30
rect 7260 0 7290 30
rect 7320 0 7350 30
rect 7380 0 7410 30
rect 7440 0 7470 30
rect 7500 0 7530 30
rect 7560 0 7590 30
rect 7620 0 7650 30
rect 7680 0 7710 30
rect 7740 0 7770 30
rect 7800 0 7830 30
rect 7860 0 7890 30
rect 7920 0 7950 30
rect 7980 0 8010 30
rect 8040 0 8070 30
rect 8100 0 8130 30
rect 8160 0 8190 30
rect 8220 0 8250 30
rect 8280 0 8310 30
rect 8340 0 8370 30
rect 8400 0 8430 30
rect 8460 0 8490 30
rect 8520 0 8550 30
rect 8580 0 8610 30
rect 8640 0 8670 30
rect 8700 0 8730 30
rect 8760 0 8790 30
rect 8820 0 8850 30
rect 8880 0 8910 30
rect 8940 0 8970 30
rect 9000 0 9030 30
rect 9060 0 9090 30
rect 9120 0 9150 30
rect 9180 0 9210 30
rect 9240 0 9270 30
rect 9300 0 9330 30
rect 9360 0 9390 30
rect 9420 0 9450 30
rect 9480 0 9510 30
rect 9540 0 9570 30
rect 9600 0 9630 30
rect 9660 0 9690 30
rect 9720 0 9750 30
rect 9780 0 9810 30
rect 9840 0 9870 30
rect 9900 0 9930 30
rect 9960 0 9990 30
rect 10020 0 10050 30
rect 10080 0 10110 30
rect 10140 0 10170 30
rect 10200 0 10230 30
rect 10260 0 10290 30
rect 10320 0 10350 30
rect 10380 0 10410 30
rect 10440 0 10470 30
rect 10500 0 10530 30
rect 10560 0 10590 30
rect 10620 0 10650 30
rect 10680 0 10730 30
use ring_osc  ring_osc_0
timestamp 1637231857
transform 1 0 300 0 1 111
box -300 -31 10550 3469
<< end >>
