magic
tech sky130A
magscale 1 2
timestamp 1623563441
<< locali >>
rect 0 20 22 80
rect 82 20 120 80
rect 180 20 220 80
rect 280 20 318 80
rect 378 20 400 80
<< viali >>
rect 22 20 82 80
rect 120 20 180 80
rect 220 20 280 80
rect 318 20 378 80
<< metal1 >>
rect 16 80 384 98
rect 16 20 22 80
rect 86 20 98 80
rect 302 20 314 80
rect 378 20 384 80
rect 16 2 384 20
<< via1 >>
rect 26 20 82 80
rect 82 20 86 80
rect 98 20 120 80
rect 120 20 158 80
rect 170 20 180 80
rect 180 20 220 80
rect 220 20 230 80
rect 242 20 280 80
rect 280 20 302 80
rect 314 20 318 80
rect 318 20 374 80
<< metal2 >>
rect 0 82 400 98
rect 0 80 36 82
rect 100 80 124 82
rect 188 80 212 82
rect 276 80 300 82
rect 364 80 400 82
rect 0 20 26 80
rect 374 20 400 80
rect 0 18 36 20
rect 100 18 124 20
rect 188 18 212 20
rect 276 18 300 20
rect 364 18 400 20
rect 0 2 400 18
<< via2 >>
rect 36 80 100 82
rect 124 80 188 82
rect 212 80 276 82
rect 300 80 364 82
rect 36 20 86 80
rect 86 20 98 80
rect 98 20 100 80
rect 124 20 158 80
rect 158 20 170 80
rect 170 20 188 80
rect 212 20 230 80
rect 230 20 242 80
rect 242 20 276 80
rect 300 20 302 80
rect 302 20 314 80
rect 314 20 364 80
rect 36 18 100 20
rect 124 18 188 20
rect 212 18 276 20
rect 300 18 364 20
<< metal3 >>
rect 0 87 400 98
rect 0 14 32 87
rect 104 14 120 87
rect 192 14 208 87
rect 280 14 296 87
rect 368 14 400 87
rect 0 2 400 14
<< via3 >>
rect 32 82 104 87
rect 32 18 36 82
rect 36 18 100 82
rect 100 18 104 82
rect 32 14 104 18
rect 120 82 192 87
rect 120 18 124 82
rect 124 18 188 82
rect 188 18 192 82
rect 120 14 192 18
rect 208 82 280 87
rect 208 18 212 82
rect 212 18 276 82
rect 276 18 280 82
rect 208 14 280 18
rect 296 82 368 87
rect 296 18 300 82
rect 300 18 364 82
rect 364 18 368 82
rect 296 14 368 18
<< metal4 >>
rect 0 87 400 98
rect 0 14 32 87
rect 104 14 120 87
rect 192 14 208 87
rect 280 14 296 87
rect 368 14 400 87
rect 0 2 400 14
<< end >>
