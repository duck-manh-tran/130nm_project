*	Cell				 	: ring oscillator testbench
*  Generated for		: NGSPICE
*  Library name		: ADC_130nm
*  Design cell name	: ring_osc_tb.spice
******************************************************

.global gnd vdd
.lib /home/LOCAL/manhtd_61d/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt 
.inc vco_w6_ext.spice
.inc sky130_digital.spice
.param mc_mm_switch=1
*_____________cross coupling inverter testbench__________________*

Xr3 p3[0] p3[1] p3[2] p3[3] p3[4] p3[5] p3[6] p3[7] p3[8] p3[9] p3[10] enb input_sig vdd gnd vco_w6_r100

X_phase_ro_0 clk p3[0] gnd vdd ro[0] phase_ro
X_phase_ro_1 clk p3[1] gnd vdd ro[1] phase_ro
X_phase_ro_2 clk p3[2] gnd vdd ro[2] phase_ro
X_phase_ro_3 clk p3[3] gnd vdd ro[3] phase_ro
X_phase_ro_4 clk p3[4] gnd vdd ro[4] phase_ro
X_phase_ro_5 clk p3[5] gnd vdd ro[5] phase_ro
X_phase_ro_6 clk p3[6] gnd vdd ro[6] phase_ro
X_phase_ro_7 clk p3[7] gnd vdd ro[7] phase_ro
X_phase_ro_8 clk p3[8] gnd vdd ro[8] phase_ro
X_phase_ro_9 clk p3[9] gnd vdd ro[9] phase_ro
X_phase_ro_10 clk p3[10] gnd vdd ro[10] phase_ro

V1 vdd gnd DC=1.8
V3 input_sig gnd SIN(0.65 0.45 11K 0 0 0)
V4 enb gnd DC=0 PULSE( 0 1.8 0 20n 20n 200n 1 )
V5 clk gnd DC=0 PULSE( 0 1.8 0 1n 1n 19n 40n )
V6 smpl_pul gnd DC=0 PULSE( 0 1.8 0 1n 1n 1n 40n )

*option INTERP
*save "ro[0]" "ro[1]" "ro[2]" "ro[3]" "ro[4]" "ro[5]" 
*+ "ro[6]" "ro[7]" "ro[8]" "ro[9]" "ro[10]" clk smpl_pul input_sig
.tran 2n 1u
*	print "ro[0]" "ro[1]" "ro[2]" > ./result/ro_vco_w6_1.txt
*	print "ro[3]" "ro[4]" "ro[5]" > ./result/ro_vco_w6_2.txt
*	print "ro[6]" "ro[7]" "ro[8]" > ./result/ro_vco_w6_3.txt
*	print "ro[9]" "ro[10]" > ./result/ro_vco_w6_4.txt
*	print clk smpl_pul > ./result/clk.txt

