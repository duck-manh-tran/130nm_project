magic
tech sky130A
magscale 1 2
timestamp 1623147612
<< nwell >>
rect -196 -220 1014 1155
<< pmos >>
rect 0 -1 380 999
rect 438 -1 818 999
<< pdiff >>
rect -58 965 0 999
rect -58 925 -46 965
rect -12 925 0 965
rect -58 891 0 925
rect -58 851 -46 891
rect -12 851 0 891
rect -58 817 0 851
rect -58 777 -46 817
rect -12 777 0 817
rect -58 743 0 777
rect -58 703 -46 743
rect -12 703 0 743
rect -58 669 0 703
rect -58 629 -46 669
rect -12 629 0 669
rect -58 595 0 629
rect -58 555 -46 595
rect -12 555 0 595
rect -58 521 0 555
rect -58 481 -46 521
rect -12 481 0 521
rect -58 447 0 481
rect -58 407 -46 447
rect -12 407 0 447
rect -58 373 0 407
rect -58 333 -46 373
rect -12 333 0 373
rect -58 299 0 333
rect -58 259 -46 299
rect -12 259 0 299
rect -58 225 0 259
rect -58 185 -46 225
rect -12 185 0 225
rect -58 151 0 185
rect -58 111 -46 151
rect -12 111 0 151
rect -58 77 0 111
rect -58 37 -46 77
rect -12 37 0 77
rect -58 -1 0 37
rect 380 965 438 999
rect 380 925 392 965
rect 426 925 438 965
rect 380 891 438 925
rect 380 851 392 891
rect 426 851 438 891
rect 380 817 438 851
rect 380 777 392 817
rect 426 777 438 817
rect 380 743 438 777
rect 380 703 392 743
rect 426 703 438 743
rect 380 669 438 703
rect 380 629 392 669
rect 426 629 438 669
rect 380 595 438 629
rect 380 555 392 595
rect 426 555 438 595
rect 380 521 438 555
rect 380 481 392 521
rect 426 481 438 521
rect 380 447 438 481
rect 380 407 392 447
rect 426 407 438 447
rect 380 373 438 407
rect 380 333 392 373
rect 426 333 438 373
rect 380 299 438 333
rect 380 259 392 299
rect 426 259 438 299
rect 380 225 438 259
rect 380 185 392 225
rect 426 185 438 225
rect 380 151 438 185
rect 380 111 392 151
rect 426 111 438 151
rect 380 77 438 111
rect 380 37 392 77
rect 426 37 438 77
rect 380 -1 438 37
rect 818 965 876 999
rect 818 925 830 965
rect 864 925 876 965
rect 818 891 876 925
rect 818 851 830 891
rect 864 851 876 891
rect 818 817 876 851
rect 818 777 830 817
rect 864 777 876 817
rect 818 743 876 777
rect 818 703 830 743
rect 864 703 876 743
rect 818 669 876 703
rect 818 629 830 669
rect 864 629 876 669
rect 818 595 876 629
rect 818 555 830 595
rect 864 555 876 595
rect 818 521 876 555
rect 818 481 830 521
rect 864 481 876 521
rect 818 447 876 481
rect 818 407 830 447
rect 864 407 876 447
rect 818 373 876 407
rect 818 333 830 373
rect 864 333 876 373
rect 818 299 876 333
rect 818 259 830 299
rect 864 259 876 299
rect 818 225 876 259
rect 818 185 830 225
rect 864 185 876 225
rect 818 151 876 185
rect 818 111 830 151
rect 864 111 876 151
rect 818 77 876 111
rect 818 37 830 77
rect 864 37 876 77
rect 818 -1 876 37
<< pdiffc >>
rect -46 925 -12 965
rect -46 851 -12 891
rect -46 777 -12 817
rect -46 703 -12 743
rect -46 629 -12 669
rect -46 555 -12 595
rect -46 481 -12 521
rect -46 407 -12 447
rect -46 333 -12 373
rect -46 259 -12 299
rect -46 185 -12 225
rect -46 111 -12 151
rect -46 37 -12 77
rect 392 925 426 965
rect 392 851 426 891
rect 392 777 426 817
rect 392 703 426 743
rect 392 629 426 669
rect 392 555 426 595
rect 392 481 426 521
rect 392 407 426 447
rect 392 333 426 373
rect 392 259 426 299
rect 392 185 426 225
rect 392 111 426 151
rect 392 37 426 77
rect 830 925 864 965
rect 830 851 864 891
rect 830 777 864 817
rect 830 703 864 743
rect 830 629 864 669
rect 830 555 864 595
rect 830 481 864 521
rect 830 407 864 447
rect 830 333 864 373
rect 830 259 864 299
rect 830 185 864 225
rect 830 111 864 151
rect 830 37 864 77
<< nsubdiff >>
rect -160 1085 -60 1119
rect -20 1085 20 1119
rect 60 1085 100 1119
rect 140 1085 180 1119
rect 220 1085 260 1119
rect 300 1085 340 1119
rect 380 1085 420 1119
rect 460 1085 500 1119
rect 540 1085 580 1119
rect 620 1085 660 1119
rect 700 1085 740 1119
rect 780 1085 820 1119
rect 860 1085 978 1119
rect -160 1039 -126 1085
rect 944 1039 978 1085
rect -160 959 -126 999
rect -160 879 -126 919
rect -160 799 -126 839
rect -160 719 -126 759
rect -160 639 -126 679
rect -160 559 -126 599
rect -160 479 -126 519
rect -160 399 -126 439
rect -160 319 -126 359
rect -160 239 -126 279
rect -160 159 -126 199
rect -160 79 -126 119
rect 944 959 978 999
rect 944 879 978 919
rect 944 799 978 839
rect 944 719 978 759
rect 944 639 978 679
rect 944 559 978 599
rect 944 479 978 519
rect 944 399 978 439
rect 944 319 978 359
rect 944 239 978 279
rect 944 159 978 199
rect 944 79 978 119
<< nsubdiffcont >>
rect -60 1085 -20 1119
rect 20 1085 60 1119
rect 100 1085 140 1119
rect 180 1085 220 1119
rect 260 1085 300 1119
rect 340 1085 380 1119
rect 420 1085 460 1119
rect 500 1085 540 1119
rect 580 1085 620 1119
rect 660 1085 700 1119
rect 740 1085 780 1119
rect 820 1085 860 1119
rect -160 999 -126 1039
rect 944 999 978 1039
rect -160 919 -126 959
rect -160 839 -126 879
rect -160 759 -126 799
rect -160 679 -126 719
rect -160 599 -126 639
rect -160 519 -126 559
rect -160 439 -126 479
rect -160 359 -126 399
rect -160 279 -126 319
rect -160 199 -126 239
rect -160 119 -126 159
rect 944 919 978 959
rect 944 839 978 879
rect 944 759 978 799
rect 944 679 978 719
rect 944 599 978 639
rect 944 519 978 559
rect 944 439 978 479
rect 944 359 978 399
rect 944 279 978 319
rect 944 199 978 239
rect 944 119 978 159
<< poly >>
rect 0 999 380 1025
rect 438 999 818 1025
rect 0 -98 380 -1
rect 438 -98 818 -1
<< locali >>
rect -160 1085 -60 1119
rect -20 1085 20 1119
rect 60 1085 100 1119
rect 140 1085 180 1119
rect 220 1085 260 1119
rect 300 1085 340 1119
rect 380 1085 420 1119
rect 460 1085 500 1119
rect 540 1085 580 1119
rect 620 1085 660 1119
rect 700 1085 740 1119
rect 780 1085 820 1119
rect 860 1085 978 1119
rect -160 1039 -126 1085
rect -160 959 -126 999
rect -160 879 -126 919
rect -160 799 -126 839
rect -160 719 -126 759
rect -160 639 -126 679
rect -160 559 -126 599
rect -160 479 -126 519
rect -160 399 -126 439
rect -160 319 -126 359
rect -160 239 -126 279
rect -160 159 -126 199
rect -160 79 -126 119
rect -58 965 0 1085
rect -58 925 -46 965
rect -12 925 0 965
rect -58 891 0 925
rect -58 851 -46 891
rect -12 851 0 891
rect -58 817 0 851
rect -58 777 -46 817
rect -12 777 0 817
rect -58 743 0 777
rect -58 703 -46 743
rect -12 703 0 743
rect -58 669 0 703
rect -58 629 -46 669
rect -12 629 0 669
rect -58 595 0 629
rect -58 555 -46 595
rect -12 555 0 595
rect -58 521 0 555
rect -58 481 -46 521
rect -12 481 0 521
rect -58 447 0 481
rect -58 407 -46 447
rect -12 407 0 447
rect -58 373 0 407
rect -58 333 -46 373
rect -12 333 0 373
rect -58 299 0 333
rect -58 259 -46 299
rect -12 259 0 299
rect -58 225 0 259
rect -58 185 -46 225
rect -12 185 0 225
rect -58 151 0 185
rect -58 111 -46 151
rect -12 111 0 151
rect -58 77 0 111
rect -58 37 -46 77
rect -12 37 0 77
rect -58 -5 0 37
rect 392 965 426 1003
rect 392 891 426 925
rect 392 817 426 851
rect 392 743 426 777
rect 392 669 426 703
rect 392 595 426 629
rect 392 521 426 555
rect 392 447 426 481
rect 392 373 426 407
rect 392 299 426 333
rect 392 225 426 259
rect 392 151 426 185
rect 392 77 426 111
rect 392 -5 426 37
rect 818 965 876 1085
rect 818 925 830 965
rect 864 925 876 965
rect 818 891 876 925
rect 818 851 830 891
rect 864 851 876 891
rect 818 817 876 851
rect 818 777 830 817
rect 864 777 876 817
rect 818 743 876 777
rect 818 703 830 743
rect 864 703 876 743
rect 818 669 876 703
rect 818 629 830 669
rect 864 629 876 669
rect 818 595 876 629
rect 818 555 830 595
rect 864 555 876 595
rect 818 521 876 555
rect 818 481 830 521
rect 864 481 876 521
rect 818 447 876 481
rect 818 407 830 447
rect 864 407 876 447
rect 818 373 876 407
rect 818 333 830 373
rect 864 333 876 373
rect 818 299 876 333
rect 818 259 830 299
rect 864 259 876 299
rect 818 225 876 259
rect 818 185 830 225
rect 864 185 876 225
rect 818 151 876 185
rect 818 111 830 151
rect 864 111 876 151
rect 818 77 876 111
rect 944 1039 978 1085
rect 944 959 978 999
rect 944 879 978 919
rect 944 799 978 839
rect 944 719 978 759
rect 944 639 978 679
rect 944 559 978 599
rect 944 479 978 519
rect 944 399 978 439
rect 944 319 978 359
rect 944 239 978 279
rect 944 159 978 199
rect 944 79 978 119
rect 818 37 830 77
rect 864 37 876 77
rect 818 -5 876 37
<< end >>
