*	Cell				 	: ring oscillator testbench
*  Generated for		: NGSPICE
*  Library name		: ADC_130nm
*  Design cell name	: ring_osc_tb.spice
******************************************************

.lib /home/dkit/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt 

.global gnd vdd
.inc sky130_digital.spice
.inc adc_130nm.spice
.param mc_mm_switch=1

*_____________cross coupling inverter testbench__________________*

Xr1 p1[0] p1[1] p1[2] p1[3] p1[4] p1[5] p1[6] p1[7] p1[8] p1[9] p1[10] input_1 enb vdd gnd vco
Xr2 p2[0] p2[1] p2[2] p2[3] p2[4] p2[5] p2[6] p2[7] p2[8] p2[9] p2[10] input_2 enb vdd gnd v_crt_v2 vco_r100
Xr3 p3[0] p3[1] p3[2] p3[3] p3[4] p3[5] p3[6] p3[7] p3[8] p3[9] p3[10] input_2 enb vdd gnd v_crt_v3 vco_w6_r100

V1 vdd gnd DC=1.8
V2 input_1 gnd DC=0.8
V3 input_2 gnd DC=0.8
V4 enb gnd DC=0 PULSE( 0 1.8 0 20n 20n 200n 1 )

.tran 0.4n 5u

.control
set num_threads=12
let prd=1
let Vin=unitvec(60)
let Vin[0]=0.1
let freq_v1=unitvec(60)
let Vcrt_v1=unitvec(60)
let freq_v2=unitvec(60)
let Vcrt_v2=unitvec(60)
let freq_v3=unitvec(60)
let Vcrt_v3=unitvec(60)
let ix=0
while Vin[ix] < 1.21
	let Vcrt_v1[ix]=Vin[ix]/2
	alter V2 DC=Vcrt_v1[ix]
	alter V3 DC=Vin[ix]
	run		
	MEAS TRAN prd TRIG p1[0] VAL=0.9 RISE=8 TARG p1[0] VAL=0.9 RISE =9
	let freq_v1[ix] = 1/prd	

	MEAS TRAN prd TRIG p2[0] VAL=0.9 RISE=8 TARG p2[0] VAL=0.9 RISE =9
	MEAS TRAN Vcrt_v2[ix] AVG v(v_crt_v2) from=3u to=4u
	let freq_v2[ix] = 1/prd

	MEAS TRAN prd TRIG p3[0] VAL=0.9 RISE=8 TARG p3[0] VAL=0.9 RISE =9
	MEAS TRAN Vcrt_v3[ix] AVG v(v_crt_v3) from=3u to=4u
	let freq_v3[ix] = 1/prd
	
	let ix = ix+1
	Let Vin[ix] = Vin[ix-1]+0.5
end

print Vin Vcrt_v1 freq_v1 > ./result/vco_test.txt
print Vin Vcrt_v2 freq_v2 > ./result/vco_r100_test.txt
print Vin Vcrt_v3 freq_v3 > ./result/vco_w6_r100_test.txt
.endc

