magic
tech sky130A
magscale 1 2
timestamp 1623529308
<< psubdiff >>
rect -20 0 60 60
rect 120 0 180 60
rect 240 0 300 60
rect 360 0 420 60
rect 480 0 540 60
rect 600 0 660 60
rect 720 0 780 60
rect 840 0 900 60
rect 960 0 1020 60
rect 1080 0 1140 60
rect 1200 0 1260 60
rect 1320 0 1380 60
rect 1440 0 1500 60
rect 1560 0 1620 60
rect 1680 0 1740 60
rect 1800 0 1860 60
rect 1920 0 1980 60
rect 2040 0 2100 60
rect 2160 0 2220 60
rect 2280 0 2340 60
rect 2400 0 2460 60
rect 2520 0 2580 60
rect 2640 0 2700 60
rect 2760 0 2820 60
rect 2880 0 2940 60
rect 3000 0 3060 60
rect 3120 0 3180 60
rect 3240 0 3300 60
rect 3360 0 3420 60
rect 3480 0 3540 60
rect 3600 0 3660 60
rect 3720 0 3780 60
rect 3840 0 3900 60
rect 3960 0 4020 60
rect 4080 0 4140 60
rect 4200 0 4260 60
rect 4320 0 4380 60
rect 4440 0 4500 60
rect 4560 0 4620 60
rect 4680 0 4740 60
rect 4800 0 4860 60
rect 4920 0 4980 60
rect 5040 0 5100 60
rect 5160 0 5220 60
rect 5280 0 5340 60
rect 5400 0 5460 60
rect 5520 0 5580 60
rect 5640 0 5700 60
rect 5760 0 5820 60
rect 5880 0 5940 60
rect 6000 0 6060 60
rect 6120 0 6180 60
rect 6240 0 6300 60
rect 6360 0 6420 60
rect 6480 0 6540 60
rect 6600 0 6660 60
rect 6720 0 6780 60
rect 6840 0 6900 60
rect 6960 0 7020 60
rect 7080 0 7140 60
rect 7200 0 7260 60
rect 7320 0 7380 60
rect 7440 0 7500 60
rect 7560 0 7620 60
rect 7680 0 7740 60
rect 7800 0 7860 60
rect 7920 0 7980 60
rect 8040 0 8100 60
rect 8160 0 8220 60
rect 8280 0 8340 60
rect 8400 0 8460 60
rect 8520 0 8580 60
rect 8640 0 8700 60
rect 8760 0 8820 60
rect 8880 0 8940 60
rect 9000 0 9060 60
rect 9120 0 9180 60
rect 9240 0 9300 60
rect 9360 0 9420 60
rect 9480 0 9540 60
rect 9600 0 9660 60
rect 9720 0 9780 60
rect 9840 0 9900 60
rect 9960 0 10020 60
rect 10080 0 10140 60
rect 10200 0 10260 60
rect 10320 0 10380 60
rect 10440 0 10500 60
rect 10560 0 10620 60
rect 10680 0 10740 60
rect 10800 0 10860 60
rect 10920 0 10980 60
rect 11040 0 11100 60
rect 11160 0 11220 60
rect 11280 0 11340 60
rect 11400 0 11460 60
rect 11520 0 11580 60
rect 11640 0 11700 60
rect 11760 0 11820 60
rect 11880 0 11940 60
rect 12000 0 12060 60
rect 12120 0 12180 60
rect 12240 0 12300 60
rect 12360 0 12420 60
rect 12480 0 12540 60
rect 12600 0 12660 60
rect 12720 0 12780 60
rect 12840 0 12900 60
rect 12960 0 13020 60
rect 13080 0 13140 60
rect 13200 0 13260 60
rect 13320 0 13380 60
rect 13440 0 13500 60
rect 13560 0 13620 60
rect 13680 0 13740 60
rect 13800 0 13860 60
rect 13920 0 13980 60
rect 14040 0 14100 60
rect 14160 0 14220 60
rect 14280 0 14340 60
rect 14400 0 14460 60
rect 14520 0 14580 60
rect 14640 0 14700 60
rect 14760 0 14820 60
rect 14880 0 14940 60
rect 15000 0 15060 60
rect 15120 0 15180 60
rect 15240 0 15300 60
rect 15360 0 15420 60
rect 15480 0 15540 60
rect 15600 0 15660 60
rect 15720 0 15780 60
rect 15840 0 15900 60
rect 15960 0 16020 60
rect 16080 0 16140 60
rect 16200 0 16260 60
rect 16320 0 16380 60
rect 16440 0 16500 60
rect 16560 0 16620 60
rect 16680 0 16740 60
rect 16800 0 16860 60
rect 16920 0 16980 60
rect 17040 0 17100 60
rect 17160 0 17220 60
rect 17280 0 17340 60
rect 17400 0 17460 60
rect 17520 0 17580 60
rect 17640 0 17700 60
rect 17760 0 17820 60
rect 17880 0 17940 60
rect 18000 0 18060 60
rect -20 -40 40 0
rect -20 -160 40 -100
rect -20 -280 40 -220
rect -20 -400 40 -340
rect -20 -520 40 -460
rect -20 -640 40 -580
rect -20 -760 40 -700
rect -20 -880 40 -820
rect -20 -1000 40 -940
rect -20 -1120 40 -1060
rect -20 -1240 40 -1180
rect -20 -1360 40 -1300
rect -20 -1480 40 -1420
rect -20 -1600 40 -1540
rect -20 -1720 40 -1660
rect -20 -1840 40 -1780
rect -20 -1960 40 -1900
rect -20 -2080 40 -2020
rect -20 -2200 40 -2140
rect -20 -2320 40 -2260
rect -20 -2440 40 -2380
rect -20 -2560 40 -2500
rect -20 -2680 40 -2620
rect -20 -2800 40 -2740
rect -20 -2920 40 -2860
rect -20 -3020 40 -2980
rect -1680 -3186 -1640 -3126
rect -1580 -3186 -1520 -3126
rect -1460 -3186 -1400 -3126
rect -1340 -3186 -1280 -3126
rect -1220 -3186 -1160 -3126
rect -1100 -3186 -1040 -3126
rect -980 -3186 -920 -3126
rect -860 -3186 -800 -3126
rect -740 -3186 -680 -3126
rect -620 -3186 -560 -3126
rect -500 -3186 -440 -3126
rect -380 -3186 -320 -3126
rect -260 -3186 -200 -3126
rect -140 -3186 -80 -3126
rect -20 -3186 40 -3080
rect 18120 -40 18180 60
rect 18120 -160 18180 -100
rect 18120 -280 18180 -220
rect 18120 -400 18180 -340
rect 18120 -520 18180 -460
rect 18120 -640 18180 -580
rect 18120 -760 18180 -700
rect 18120 -880 18180 -820
rect 18120 -1000 18180 -940
rect 18120 -1120 18180 -1060
rect 18120 -1240 18180 -1180
rect 18120 -1360 18180 -1300
rect 18120 -1480 18180 -1420
rect 18120 -1600 18180 -1540
rect 18120 -1720 18180 -1660
rect 18120 -1840 18180 -1780
rect 18120 -1960 18180 -1900
rect 18120 -2080 18180 -2020
rect 18120 -2200 18180 -2140
rect 18120 -2320 18180 -2260
rect 18120 -2440 18180 -2380
rect 18120 -2560 18180 -2500
rect 18120 -2680 18180 -2620
rect 18120 -2800 18180 -2740
rect 18120 -2920 18180 -2860
rect 18120 -3020 18180 -2980
rect 18120 -3126 18180 -3080
rect 100 -3186 140 -3126
rect 200 -3186 260 -3126
rect 320 -3186 380 -3126
rect 440 -3186 500 -3126
rect 560 -3186 620 -3126
rect 680 -3186 740 -3126
rect 800 -3186 860 -3126
rect 920 -3186 980 -3126
rect 1040 -3186 1100 -3126
rect 1160 -3186 1220 -3126
rect 1280 -3186 1340 -3126
rect 1400 -3186 1460 -3126
rect 1520 -3186 1580 -3126
rect 1640 -3186 1700 -3126
rect 1760 -3186 1820 -3126
rect 1880 -3186 1940 -3126
rect 2000 -3186 2060 -3126
rect 2120 -3186 2180 -3126
rect 2240 -3186 2300 -3126
rect 2360 -3186 2420 -3126
rect 2480 -3186 2540 -3126
rect 2600 -3186 2660 -3126
rect 2720 -3186 2780 -3126
rect 2840 -3186 2900 -3126
rect 2960 -3186 3020 -3126
rect 3080 -3186 3140 -3126
rect 3200 -3186 3260 -3126
rect 3320 -3186 3380 -3126
rect 3440 -3186 3500 -3126
rect 3560 -3186 3620 -3126
rect 3680 -3186 3740 -3126
rect 3800 -3186 3860 -3126
rect 3920 -3186 3980 -3126
rect 4040 -3186 4100 -3126
rect 4160 -3186 4220 -3126
rect 4280 -3186 4340 -3126
rect 4400 -3186 4460 -3126
rect 4520 -3186 4580 -3126
rect 4640 -3186 4700 -3126
rect 4760 -3186 4820 -3126
rect 4880 -3186 4940 -3126
rect 5000 -3186 5060 -3126
rect 5120 -3186 5180 -3126
rect 5240 -3186 5300 -3126
rect 5360 -3186 5420 -3126
rect 5480 -3186 5540 -3126
rect 5600 -3186 5660 -3126
rect 5720 -3186 5780 -3126
rect 5840 -3186 5900 -3126
rect 5960 -3186 6020 -3126
rect 6080 -3186 6140 -3126
rect 6200 -3186 6260 -3126
rect 6320 -3186 6380 -3126
rect 6440 -3186 6500 -3126
rect 6560 -3186 6620 -3126
rect 6680 -3186 6740 -3126
rect 6800 -3186 6860 -3126
rect 6920 -3186 6980 -3126
rect 7040 -3186 7100 -3126
rect 7160 -3186 7220 -3126
rect 7280 -3186 7340 -3126
rect 7400 -3186 7460 -3126
rect 7520 -3186 7580 -3126
rect 7640 -3186 7700 -3126
rect 7760 -3186 7820 -3126
rect 7880 -3186 7940 -3126
rect 8000 -3186 8060 -3126
rect 8120 -3186 8180 -3126
rect 8240 -3186 8300 -3126
rect 8360 -3186 8420 -3126
rect 8480 -3186 8540 -3126
rect 8600 -3186 8660 -3126
rect 8720 -3186 8780 -3126
rect 8840 -3186 8900 -3126
rect 8960 -3186 9020 -3126
rect 9080 -3186 9140 -3126
rect 9200 -3186 9260 -3126
rect 9320 -3186 9380 -3126
rect 9440 -3186 9500 -3126
rect 9560 -3186 9620 -3126
rect 9680 -3186 9740 -3126
rect 9800 -3186 9860 -3126
rect 9920 -3186 9980 -3126
rect 10040 -3186 10100 -3126
rect 10160 -3186 10220 -3126
rect 10280 -3186 10340 -3126
rect 10400 -3186 10460 -3126
rect 10520 -3186 10580 -3126
rect 10640 -3186 10700 -3126
rect 10760 -3186 10820 -3126
rect 10880 -3186 10940 -3126
rect 11000 -3186 11060 -3126
rect 11120 -3186 11180 -3126
rect 11240 -3186 11300 -3126
rect 11360 -3186 11420 -3126
rect 11480 -3186 11540 -3126
rect 11600 -3186 11660 -3126
rect 11720 -3186 11780 -3126
rect 11840 -3186 11900 -3126
rect 11960 -3186 12020 -3126
rect 12080 -3186 12140 -3126
rect 12200 -3186 12260 -3126
rect 12320 -3186 12380 -3126
rect 12440 -3186 12500 -3126
rect 12560 -3186 12620 -3126
rect 12680 -3186 12740 -3126
rect 12800 -3186 12860 -3126
rect 12920 -3186 12980 -3126
rect 13040 -3186 13100 -3126
rect 13160 -3186 13220 -3126
rect 13280 -3186 13340 -3126
rect 13400 -3186 13460 -3126
rect 13520 -3186 13580 -3126
rect 13640 -3186 13700 -3126
rect 13760 -3186 13820 -3126
rect 13880 -3186 13940 -3126
rect 14000 -3186 14060 -3126
rect 14120 -3186 14180 -3126
rect 14240 -3186 14300 -3126
rect 14360 -3186 14420 -3126
rect 14480 -3186 14540 -3126
rect 14600 -3186 14660 -3126
rect 14720 -3186 14780 -3126
rect 14840 -3186 14900 -3126
rect 14960 -3186 15020 -3126
rect 15080 -3186 15140 -3126
rect 15200 -3186 15260 -3126
rect 15320 -3186 15380 -3126
rect 15440 -3186 15500 -3126
rect 15560 -3186 15620 -3126
rect 15680 -3186 15740 -3126
rect 15800 -3186 15860 -3126
rect 15920 -3186 15980 -3126
rect 16040 -3186 16100 -3126
rect 16160 -3186 16220 -3126
rect 16280 -3186 16340 -3126
rect 16400 -3186 16460 -3126
rect 16520 -3186 16580 -3126
rect 16640 -3186 16700 -3126
rect 16760 -3186 16820 -3126
rect 16880 -3186 16940 -3126
rect 17000 -3186 17060 -3126
rect 17120 -3186 17180 -3126
rect 17240 -3186 17300 -3126
rect 17360 -3186 17420 -3126
rect 17480 -3186 17540 -3126
rect 17600 -3186 17660 -3126
rect 17720 -3186 17780 -3126
rect 17840 -3186 17900 -3126
rect 17960 -3186 18020 -3126
rect 18080 -3186 18140 -3126
rect 18200 -3186 18260 -3126
rect 18320 -3186 18380 -3126
rect 18440 -3186 18500 -3126
rect 18560 -3186 18620 -3126
rect 18680 -3186 18740 -3126
rect 18800 -3186 18860 -3126
rect 18920 -3186 18980 -3126
rect 19040 -3186 19100 -3126
rect 19160 -3186 19220 -3126
rect 19280 -3186 19340 -3126
rect 19400 -3186 19460 -3126
rect 19520 -3186 19580 -3126
rect 19640 -3186 19700 -3126
rect 19760 -3186 19820 -3126
rect 19880 -3186 19940 -3126
rect 20000 -3186 20060 -3126
rect 20120 -3186 20145 -3126
rect -1680 -3226 -1620 -3186
rect -1680 -3346 -1620 -3286
rect -1680 -3466 -1620 -3406
rect -1680 -3586 -1620 -3526
rect -1680 -3706 -1620 -3646
rect -1680 -3826 -1620 -3766
rect -1680 -3946 -1620 -3886
rect -1680 -4066 -1620 -4006
rect -1680 -4186 -1620 -4126
rect -1680 -4306 -1620 -4246
rect -1680 -4426 -1620 -4366
rect -1680 -4546 -1620 -4486
rect -1680 -4666 -1620 -4606
rect -1680 -4786 -1620 -4726
rect -1680 -4906 -1620 -4846
rect -1680 -5026 -1620 -4966
rect -1680 -5146 -1620 -5086
rect -1680 -5266 -1620 -5206
rect -1680 -5386 -1620 -5326
rect -1680 -5506 -1620 -5446
rect -1680 -5626 -1620 -5566
rect -1680 -5746 -1620 -5686
rect -1680 -5866 -1620 -5806
rect -1680 -5986 -1620 -5926
rect -1680 -6106 -1620 -6046
rect -1680 -6206 -1620 -6166
rect -1680 -6360 -1620 -6266
rect 20080 -3200 20145 -3186
rect 20080 -3246 20140 -3200
rect 20080 -3366 20140 -3306
rect 20080 -3486 20140 -3426
rect 20080 -3606 20140 -3546
rect 20080 -3726 20140 -3666
rect 20080 -3846 20140 -3786
rect 20080 -3966 20140 -3906
rect 20080 -4086 20140 -4026
rect 20080 -4206 20140 -4146
rect 20080 -4326 20140 -4266
rect 20080 -4446 20140 -4386
rect 20080 -4566 20140 -4506
rect 20080 -4686 20140 -4626
rect 20080 -4806 20140 -4746
rect 20080 -4926 20140 -4866
rect 20080 -5046 20140 -4986
rect 20080 -5166 20140 -5106
rect 20080 -5286 20140 -5226
rect 20080 -5406 20140 -5346
rect 20080 -5526 20140 -5466
rect 20080 -5646 20140 -5586
rect 20080 -5766 20140 -5706
rect 20080 -5886 20140 -5826
rect 20080 -6006 20140 -5946
rect 20080 -6126 20140 -6066
rect 20080 -6240 20140 -6186
rect -1560 -6360 -1500 -6300
rect -1440 -6360 -1380 -6300
rect -1320 -6360 -1260 -6300
rect -1200 -6360 -1140 -6300
rect -1080 -6360 -1020 -6300
rect -960 -6360 -900 -6300
rect -840 -6360 -780 -6300
rect -720 -6360 -660 -6300
rect -600 -6360 -540 -6300
rect -480 -6360 -420 -6300
rect -360 -6360 -300 -6300
rect -240 -6360 -180 -6300
rect -120 -6360 -60 -6300
rect 0 -6360 60 -6300
rect 120 -6360 180 -6300
rect 240 -6360 300 -6300
rect 360 -6360 420 -6300
rect 480 -6360 540 -6300
rect 600 -6360 660 -6300
rect 720 -6360 780 -6300
rect 840 -6360 900 -6300
rect 960 -6360 1020 -6300
rect 1080 -6360 1140 -6300
rect 1200 -6360 1260 -6300
rect 1320 -6360 1380 -6300
rect 1440 -6360 1500 -6300
rect 1560 -6360 1620 -6300
rect 1680 -6360 1740 -6300
rect 1800 -6360 1860 -6300
rect 1920 -6360 1980 -6300
rect 2040 -6360 2100 -6300
rect 2160 -6360 2220 -6300
rect 2280 -6360 2340 -6300
rect 2400 -6360 2460 -6300
rect 2520 -6360 2580 -6300
rect 2640 -6360 2700 -6300
rect 2760 -6360 2820 -6300
rect 2880 -6360 2940 -6300
rect 3000 -6360 3060 -6300
rect 3120 -6360 3180 -6300
rect 3240 -6360 3300 -6300
rect 3360 -6360 3420 -6300
rect 3480 -6360 3540 -6300
rect 3600 -6360 3660 -6300
rect 3720 -6360 3780 -6300
rect 3840 -6360 3900 -6300
rect 3960 -6360 4020 -6300
rect 4080 -6360 4140 -6300
rect 4200 -6360 4260 -6300
rect 4320 -6360 4380 -6300
rect 4440 -6360 4500 -6300
rect 4560 -6360 4620 -6300
rect 4680 -6360 4740 -6300
rect 4800 -6360 4860 -6300
rect 4920 -6360 4980 -6300
rect 5040 -6360 5100 -6300
rect 5160 -6360 5220 -6300
rect 5280 -6360 5340 -6300
rect 5400 -6360 5460 -6300
rect 5520 -6360 5580 -6300
rect 5640 -6360 5700 -6300
rect 5760 -6360 5820 -6300
rect 5880 -6360 5940 -6300
rect 6000 -6360 6060 -6300
rect 6120 -6360 6180 -6300
rect 6240 -6360 6300 -6300
rect 6360 -6360 6420 -6300
rect 6480 -6360 6540 -6300
rect 6600 -6360 6660 -6300
rect 6720 -6360 6780 -6300
rect 6840 -6360 6900 -6300
rect 6960 -6360 7020 -6300
rect 7080 -6360 7140 -6300
rect 7200 -6360 7260 -6300
rect 7320 -6360 7380 -6300
rect 7440 -6360 7500 -6300
rect 7560 -6360 7620 -6300
rect 7680 -6360 7740 -6300
rect 7800 -6360 7860 -6300
rect 7920 -6360 7980 -6300
rect 8040 -6360 8100 -6300
rect 8160 -6360 8220 -6300
rect 8280 -6360 8340 -6300
rect 8400 -6360 8460 -6300
rect 8520 -6360 8580 -6300
rect 8640 -6360 8700 -6300
rect 8760 -6360 8820 -6300
rect 8880 -6360 8940 -6300
rect 9000 -6360 9060 -6300
rect 9120 -6360 9180 -6300
rect 9240 -6360 9300 -6300
rect 9360 -6360 9420 -6300
rect 9480 -6360 9540 -6300
rect 9600 -6360 9660 -6300
rect 9720 -6360 9780 -6300
rect 9840 -6360 9900 -6300
rect 9960 -6360 10020 -6300
rect 10080 -6360 10140 -6300
rect 10200 -6360 10260 -6300
rect 10320 -6360 10380 -6300
rect 10440 -6360 10500 -6300
rect 10560 -6360 10620 -6300
rect 10680 -6360 10740 -6300
rect 10800 -6360 10860 -6300
rect 10920 -6360 10980 -6300
rect 11040 -6360 11100 -6300
rect 11160 -6360 11220 -6300
rect 11280 -6360 11340 -6300
rect 11400 -6360 11460 -6300
rect 11520 -6360 11580 -6300
rect 11640 -6360 11700 -6300
rect 11760 -6360 11820 -6300
rect 11880 -6360 11940 -6300
rect 12000 -6360 12060 -6300
rect 12120 -6360 12180 -6300
rect 12240 -6360 12300 -6300
rect 12360 -6360 12420 -6300
rect 12480 -6360 12540 -6300
rect 12600 -6360 12660 -6300
rect 12720 -6360 12780 -6300
rect 12840 -6360 12900 -6300
rect 12960 -6360 13020 -6300
rect 13080 -6360 13140 -6300
rect 13200 -6360 13260 -6300
rect 13320 -6360 13380 -6300
rect 13440 -6360 13500 -6300
rect 13560 -6360 13620 -6300
rect 13680 -6360 13740 -6300
rect 13800 -6360 13860 -6300
rect 13920 -6360 13980 -6300
rect 14040 -6360 14100 -6300
rect 14160 -6360 14220 -6300
rect 14280 -6360 14340 -6300
rect 14400 -6360 14460 -6300
rect 14520 -6360 14580 -6300
rect 14640 -6360 14700 -6300
rect 14760 -6360 14820 -6300
rect 14880 -6360 14940 -6300
rect 15000 -6360 15060 -6300
rect 15120 -6360 15180 -6300
rect 15240 -6360 15300 -6300
rect 15360 -6360 15420 -6300
rect 15480 -6360 15540 -6300
rect 15600 -6360 15660 -6300
rect 15720 -6360 15780 -6300
rect 15840 -6360 15900 -6300
rect 15960 -6360 16020 -6300
rect 16080 -6360 16140 -6300
rect 16200 -6360 16260 -6300
rect 16320 -6360 16380 -6300
rect 16440 -6360 16500 -6300
rect 16560 -6360 16620 -6300
rect 16680 -6360 16740 -6300
rect 16800 -6360 16860 -6300
rect 16920 -6360 16980 -6300
rect 17040 -6360 17100 -6300
rect 17160 -6360 17220 -6300
rect 17280 -6360 17340 -6300
rect 17400 -6360 17460 -6300
rect 17520 -6360 17580 -6300
rect 17640 -6360 17700 -6300
rect 17760 -6360 17820 -6300
rect 17880 -6360 17940 -6300
rect 18000 -6360 18060 -6300
rect 18120 -6360 18180 -6300
rect 18240 -6360 18300 -6300
rect 18360 -6360 18420 -6300
rect 18480 -6360 18540 -6300
rect 18600 -6360 18660 -6300
rect 18720 -6360 18780 -6300
rect 18840 -6360 18900 -6300
rect 18960 -6360 19020 -6300
rect 19080 -6360 19140 -6300
rect 19200 -6360 19260 -6300
rect 19320 -6360 19380 -6300
rect 19440 -6360 19500 -6300
rect 19560 -6360 19620 -6300
rect 19680 -6360 19740 -6300
rect 19800 -6360 19860 -6300
rect 19920 -6360 19980 -6300
rect 20040 -6360 20140 -6300
<< psubdiffcont >>
rect 60 0 120 60
rect 180 0 240 60
rect 300 0 360 60
rect 420 0 480 60
rect 540 0 600 60
rect 660 0 720 60
rect 780 0 840 60
rect 900 0 960 60
rect 1020 0 1080 60
rect 1140 0 1200 60
rect 1260 0 1320 60
rect 1380 0 1440 60
rect 1500 0 1560 60
rect 1620 0 1680 60
rect 1740 0 1800 60
rect 1860 0 1920 60
rect 1980 0 2040 60
rect 2100 0 2160 60
rect 2220 0 2280 60
rect 2340 0 2400 60
rect 2460 0 2520 60
rect 2580 0 2640 60
rect 2700 0 2760 60
rect 2820 0 2880 60
rect 2940 0 3000 60
rect 3060 0 3120 60
rect 3180 0 3240 60
rect 3300 0 3360 60
rect 3420 0 3480 60
rect 3540 0 3600 60
rect 3660 0 3720 60
rect 3780 0 3840 60
rect 3900 0 3960 60
rect 4020 0 4080 60
rect 4140 0 4200 60
rect 4260 0 4320 60
rect 4380 0 4440 60
rect 4500 0 4560 60
rect 4620 0 4680 60
rect 4740 0 4800 60
rect 4860 0 4920 60
rect 4980 0 5040 60
rect 5100 0 5160 60
rect 5220 0 5280 60
rect 5340 0 5400 60
rect 5460 0 5520 60
rect 5580 0 5640 60
rect 5700 0 5760 60
rect 5820 0 5880 60
rect 5940 0 6000 60
rect 6060 0 6120 60
rect 6180 0 6240 60
rect 6300 0 6360 60
rect 6420 0 6480 60
rect 6540 0 6600 60
rect 6660 0 6720 60
rect 6780 0 6840 60
rect 6900 0 6960 60
rect 7020 0 7080 60
rect 7140 0 7200 60
rect 7260 0 7320 60
rect 7380 0 7440 60
rect 7500 0 7560 60
rect 7620 0 7680 60
rect 7740 0 7800 60
rect 7860 0 7920 60
rect 7980 0 8040 60
rect 8100 0 8160 60
rect 8220 0 8280 60
rect 8340 0 8400 60
rect 8460 0 8520 60
rect 8580 0 8640 60
rect 8700 0 8760 60
rect 8820 0 8880 60
rect 8940 0 9000 60
rect 9060 0 9120 60
rect 9180 0 9240 60
rect 9300 0 9360 60
rect 9420 0 9480 60
rect 9540 0 9600 60
rect 9660 0 9720 60
rect 9780 0 9840 60
rect 9900 0 9960 60
rect 10020 0 10080 60
rect 10140 0 10200 60
rect 10260 0 10320 60
rect 10380 0 10440 60
rect 10500 0 10560 60
rect 10620 0 10680 60
rect 10740 0 10800 60
rect 10860 0 10920 60
rect 10980 0 11040 60
rect 11100 0 11160 60
rect 11220 0 11280 60
rect 11340 0 11400 60
rect 11460 0 11520 60
rect 11580 0 11640 60
rect 11700 0 11760 60
rect 11820 0 11880 60
rect 11940 0 12000 60
rect 12060 0 12120 60
rect 12180 0 12240 60
rect 12300 0 12360 60
rect 12420 0 12480 60
rect 12540 0 12600 60
rect 12660 0 12720 60
rect 12780 0 12840 60
rect 12900 0 12960 60
rect 13020 0 13080 60
rect 13140 0 13200 60
rect 13260 0 13320 60
rect 13380 0 13440 60
rect 13500 0 13560 60
rect 13620 0 13680 60
rect 13740 0 13800 60
rect 13860 0 13920 60
rect 13980 0 14040 60
rect 14100 0 14160 60
rect 14220 0 14280 60
rect 14340 0 14400 60
rect 14460 0 14520 60
rect 14580 0 14640 60
rect 14700 0 14760 60
rect 14820 0 14880 60
rect 14940 0 15000 60
rect 15060 0 15120 60
rect 15180 0 15240 60
rect 15300 0 15360 60
rect 15420 0 15480 60
rect 15540 0 15600 60
rect 15660 0 15720 60
rect 15780 0 15840 60
rect 15900 0 15960 60
rect 16020 0 16080 60
rect 16140 0 16200 60
rect 16260 0 16320 60
rect 16380 0 16440 60
rect 16500 0 16560 60
rect 16620 0 16680 60
rect 16740 0 16800 60
rect 16860 0 16920 60
rect 16980 0 17040 60
rect 17100 0 17160 60
rect 17220 0 17280 60
rect 17340 0 17400 60
rect 17460 0 17520 60
rect 17580 0 17640 60
rect 17700 0 17760 60
rect 17820 0 17880 60
rect 17940 0 18000 60
rect 18060 0 18120 60
rect -20 -100 40 -40
rect -20 -220 40 -160
rect -20 -340 40 -280
rect -20 -460 40 -400
rect -20 -580 40 -520
rect -20 -700 40 -640
rect -20 -820 40 -760
rect -20 -940 40 -880
rect -20 -1060 40 -1000
rect -20 -1180 40 -1120
rect -20 -1300 40 -1240
rect -20 -1420 40 -1360
rect -20 -1540 40 -1480
rect -20 -1660 40 -1600
rect -20 -1780 40 -1720
rect -20 -1900 40 -1840
rect -20 -2020 40 -1960
rect -20 -2140 40 -2080
rect -20 -2260 40 -2200
rect -20 -2380 40 -2320
rect -20 -2500 40 -2440
rect -20 -2620 40 -2560
rect -20 -2740 40 -2680
rect -20 -2860 40 -2800
rect -20 -2980 40 -2920
rect -20 -3080 40 -3020
rect -1640 -3186 -1580 -3126
rect -1520 -3186 -1460 -3126
rect -1400 -3186 -1340 -3126
rect -1280 -3186 -1220 -3126
rect -1160 -3186 -1100 -3126
rect -1040 -3186 -980 -3126
rect -920 -3186 -860 -3126
rect -800 -3186 -740 -3126
rect -680 -3186 -620 -3126
rect -560 -3186 -500 -3126
rect -440 -3186 -380 -3126
rect -320 -3186 -260 -3126
rect -200 -3186 -140 -3126
rect -80 -3186 -20 -3126
rect 18120 -100 18180 -40
rect 18120 -220 18180 -160
rect 18120 -340 18180 -280
rect 18120 -460 18180 -400
rect 18120 -580 18180 -520
rect 18120 -700 18180 -640
rect 18120 -820 18180 -760
rect 18120 -940 18180 -880
rect 18120 -1060 18180 -1000
rect 18120 -1180 18180 -1120
rect 18120 -1300 18180 -1240
rect 18120 -1420 18180 -1360
rect 18120 -1540 18180 -1480
rect 18120 -1660 18180 -1600
rect 18120 -1780 18180 -1720
rect 18120 -1900 18180 -1840
rect 18120 -2020 18180 -1960
rect 18120 -2140 18180 -2080
rect 18120 -2260 18180 -2200
rect 18120 -2380 18180 -2320
rect 18120 -2500 18180 -2440
rect 18120 -2620 18180 -2560
rect 18120 -2740 18180 -2680
rect 18120 -2860 18180 -2800
rect 18120 -2980 18180 -2920
rect 18120 -3080 18180 -3020
rect 40 -3186 100 -3126
rect 140 -3186 200 -3126
rect 260 -3186 320 -3126
rect 380 -3186 440 -3126
rect 500 -3186 560 -3126
rect 620 -3186 680 -3126
rect 740 -3186 800 -3126
rect 860 -3186 920 -3126
rect 980 -3186 1040 -3126
rect 1100 -3186 1160 -3126
rect 1220 -3186 1280 -3126
rect 1340 -3186 1400 -3126
rect 1460 -3186 1520 -3126
rect 1580 -3186 1640 -3126
rect 1700 -3186 1760 -3126
rect 1820 -3186 1880 -3126
rect 1940 -3186 2000 -3126
rect 2060 -3186 2120 -3126
rect 2180 -3186 2240 -3126
rect 2300 -3186 2360 -3126
rect 2420 -3186 2480 -3126
rect 2540 -3186 2600 -3126
rect 2660 -3186 2720 -3126
rect 2780 -3186 2840 -3126
rect 2900 -3186 2960 -3126
rect 3020 -3186 3080 -3126
rect 3140 -3186 3200 -3126
rect 3260 -3186 3320 -3126
rect 3380 -3186 3440 -3126
rect 3500 -3186 3560 -3126
rect 3620 -3186 3680 -3126
rect 3740 -3186 3800 -3126
rect 3860 -3186 3920 -3126
rect 3980 -3186 4040 -3126
rect 4100 -3186 4160 -3126
rect 4220 -3186 4280 -3126
rect 4340 -3186 4400 -3126
rect 4460 -3186 4520 -3126
rect 4580 -3186 4640 -3126
rect 4700 -3186 4760 -3126
rect 4820 -3186 4880 -3126
rect 4940 -3186 5000 -3126
rect 5060 -3186 5120 -3126
rect 5180 -3186 5240 -3126
rect 5300 -3186 5360 -3126
rect 5420 -3186 5480 -3126
rect 5540 -3186 5600 -3126
rect 5660 -3186 5720 -3126
rect 5780 -3186 5840 -3126
rect 5900 -3186 5960 -3126
rect 6020 -3186 6080 -3126
rect 6140 -3186 6200 -3126
rect 6260 -3186 6320 -3126
rect 6380 -3186 6440 -3126
rect 6500 -3186 6560 -3126
rect 6620 -3186 6680 -3126
rect 6740 -3186 6800 -3126
rect 6860 -3186 6920 -3126
rect 6980 -3186 7040 -3126
rect 7100 -3186 7160 -3126
rect 7220 -3186 7280 -3126
rect 7340 -3186 7400 -3126
rect 7460 -3186 7520 -3126
rect 7580 -3186 7640 -3126
rect 7700 -3186 7760 -3126
rect 7820 -3186 7880 -3126
rect 7940 -3186 8000 -3126
rect 8060 -3186 8120 -3126
rect 8180 -3186 8240 -3126
rect 8300 -3186 8360 -3126
rect 8420 -3186 8480 -3126
rect 8540 -3186 8600 -3126
rect 8660 -3186 8720 -3126
rect 8780 -3186 8840 -3126
rect 8900 -3186 8960 -3126
rect 9020 -3186 9080 -3126
rect 9140 -3186 9200 -3126
rect 9260 -3186 9320 -3126
rect 9380 -3186 9440 -3126
rect 9500 -3186 9560 -3126
rect 9620 -3186 9680 -3126
rect 9740 -3186 9800 -3126
rect 9860 -3186 9920 -3126
rect 9980 -3186 10040 -3126
rect 10100 -3186 10160 -3126
rect 10220 -3186 10280 -3126
rect 10340 -3186 10400 -3126
rect 10460 -3186 10520 -3126
rect 10580 -3186 10640 -3126
rect 10700 -3186 10760 -3126
rect 10820 -3186 10880 -3126
rect 10940 -3186 11000 -3126
rect 11060 -3186 11120 -3126
rect 11180 -3186 11240 -3126
rect 11300 -3186 11360 -3126
rect 11420 -3186 11480 -3126
rect 11540 -3186 11600 -3126
rect 11660 -3186 11720 -3126
rect 11780 -3186 11840 -3126
rect 11900 -3186 11960 -3126
rect 12020 -3186 12080 -3126
rect 12140 -3186 12200 -3126
rect 12260 -3186 12320 -3126
rect 12380 -3186 12440 -3126
rect 12500 -3186 12560 -3126
rect 12620 -3186 12680 -3126
rect 12740 -3186 12800 -3126
rect 12860 -3186 12920 -3126
rect 12980 -3186 13040 -3126
rect 13100 -3186 13160 -3126
rect 13220 -3186 13280 -3126
rect 13340 -3186 13400 -3126
rect 13460 -3186 13520 -3126
rect 13580 -3186 13640 -3126
rect 13700 -3186 13760 -3126
rect 13820 -3186 13880 -3126
rect 13940 -3186 14000 -3126
rect 14060 -3186 14120 -3126
rect 14180 -3186 14240 -3126
rect 14300 -3186 14360 -3126
rect 14420 -3186 14480 -3126
rect 14540 -3186 14600 -3126
rect 14660 -3186 14720 -3126
rect 14780 -3186 14840 -3126
rect 14900 -3186 14960 -3126
rect 15020 -3186 15080 -3126
rect 15140 -3186 15200 -3126
rect 15260 -3186 15320 -3126
rect 15380 -3186 15440 -3126
rect 15500 -3186 15560 -3126
rect 15620 -3186 15680 -3126
rect 15740 -3186 15800 -3126
rect 15860 -3186 15920 -3126
rect 15980 -3186 16040 -3126
rect 16100 -3186 16160 -3126
rect 16220 -3186 16280 -3126
rect 16340 -3186 16400 -3126
rect 16460 -3186 16520 -3126
rect 16580 -3186 16640 -3126
rect 16700 -3186 16760 -3126
rect 16820 -3186 16880 -3126
rect 16940 -3186 17000 -3126
rect 17060 -3186 17120 -3126
rect 17180 -3186 17240 -3126
rect 17300 -3186 17360 -3126
rect 17420 -3186 17480 -3126
rect 17540 -3186 17600 -3126
rect 17660 -3186 17720 -3126
rect 17780 -3186 17840 -3126
rect 17900 -3186 17960 -3126
rect 18020 -3186 18080 -3126
rect 18140 -3186 18200 -3126
rect 18260 -3186 18320 -3126
rect 18380 -3186 18440 -3126
rect 18500 -3186 18560 -3126
rect 18620 -3186 18680 -3126
rect 18740 -3186 18800 -3126
rect 18860 -3186 18920 -3126
rect 18980 -3186 19040 -3126
rect 19100 -3186 19160 -3126
rect 19220 -3186 19280 -3126
rect 19340 -3186 19400 -3126
rect 19460 -3186 19520 -3126
rect 19580 -3186 19640 -3126
rect 19700 -3186 19760 -3126
rect 19820 -3186 19880 -3126
rect 19940 -3186 20000 -3126
rect 20060 -3186 20120 -3126
rect -1680 -3286 -1620 -3226
rect -1680 -3406 -1620 -3346
rect -1680 -3526 -1620 -3466
rect -1680 -3646 -1620 -3586
rect -1680 -3766 -1620 -3706
rect -1680 -3886 -1620 -3826
rect -1680 -4006 -1620 -3946
rect -1680 -4126 -1620 -4066
rect -1680 -4246 -1620 -4186
rect -1680 -4366 -1620 -4306
rect -1680 -4486 -1620 -4426
rect -1680 -4606 -1620 -4546
rect -1680 -4726 -1620 -4666
rect -1680 -4846 -1620 -4786
rect -1680 -4966 -1620 -4906
rect -1680 -5086 -1620 -5026
rect -1680 -5206 -1620 -5146
rect -1680 -5326 -1620 -5266
rect -1680 -5446 -1620 -5386
rect -1680 -5566 -1620 -5506
rect -1680 -5686 -1620 -5626
rect -1680 -5806 -1620 -5746
rect -1680 -5926 -1620 -5866
rect -1680 -6046 -1620 -5986
rect -1680 -6166 -1620 -6106
rect -1680 -6266 -1620 -6206
rect 20080 -3306 20140 -3246
rect 20080 -3426 20140 -3366
rect 20080 -3546 20140 -3486
rect 20080 -3666 20140 -3606
rect 20080 -3786 20140 -3726
rect 20080 -3906 20140 -3846
rect 20080 -4026 20140 -3966
rect 20080 -4146 20140 -4086
rect 20080 -4266 20140 -4206
rect 20080 -4386 20140 -4326
rect 20080 -4506 20140 -4446
rect 20080 -4626 20140 -4566
rect 20080 -4746 20140 -4686
rect 20080 -4866 20140 -4806
rect 20080 -4986 20140 -4926
rect 20080 -5106 20140 -5046
rect 20080 -5226 20140 -5166
rect 20080 -5346 20140 -5286
rect 20080 -5466 20140 -5406
rect 20080 -5586 20140 -5526
rect 20080 -5706 20140 -5646
rect 20080 -5826 20140 -5766
rect 20080 -5946 20140 -5886
rect 20080 -6066 20140 -6006
rect 20080 -6186 20140 -6126
rect 20080 -6300 20140 -6240
rect -1620 -6360 -1560 -6300
rect -1500 -6360 -1440 -6300
rect -1380 -6360 -1320 -6300
rect -1260 -6360 -1200 -6300
rect -1140 -6360 -1080 -6300
rect -1020 -6360 -960 -6300
rect -900 -6360 -840 -6300
rect -780 -6360 -720 -6300
rect -660 -6360 -600 -6300
rect -540 -6360 -480 -6300
rect -420 -6360 -360 -6300
rect -300 -6360 -240 -6300
rect -180 -6360 -120 -6300
rect -60 -6360 0 -6300
rect 60 -6360 120 -6300
rect 180 -6360 240 -6300
rect 300 -6360 360 -6300
rect 420 -6360 480 -6300
rect 540 -6360 600 -6300
rect 660 -6360 720 -6300
rect 780 -6360 840 -6300
rect 900 -6360 960 -6300
rect 1020 -6360 1080 -6300
rect 1140 -6360 1200 -6300
rect 1260 -6360 1320 -6300
rect 1380 -6360 1440 -6300
rect 1500 -6360 1560 -6300
rect 1620 -6360 1680 -6300
rect 1740 -6360 1800 -6300
rect 1860 -6360 1920 -6300
rect 1980 -6360 2040 -6300
rect 2100 -6360 2160 -6300
rect 2220 -6360 2280 -6300
rect 2340 -6360 2400 -6300
rect 2460 -6360 2520 -6300
rect 2580 -6360 2640 -6300
rect 2700 -6360 2760 -6300
rect 2820 -6360 2880 -6300
rect 2940 -6360 3000 -6300
rect 3060 -6360 3120 -6300
rect 3180 -6360 3240 -6300
rect 3300 -6360 3360 -6300
rect 3420 -6360 3480 -6300
rect 3540 -6360 3600 -6300
rect 3660 -6360 3720 -6300
rect 3780 -6360 3840 -6300
rect 3900 -6360 3960 -6300
rect 4020 -6360 4080 -6300
rect 4140 -6360 4200 -6300
rect 4260 -6360 4320 -6300
rect 4380 -6360 4440 -6300
rect 4500 -6360 4560 -6300
rect 4620 -6360 4680 -6300
rect 4740 -6360 4800 -6300
rect 4860 -6360 4920 -6300
rect 4980 -6360 5040 -6300
rect 5100 -6360 5160 -6300
rect 5220 -6360 5280 -6300
rect 5340 -6360 5400 -6300
rect 5460 -6360 5520 -6300
rect 5580 -6360 5640 -6300
rect 5700 -6360 5760 -6300
rect 5820 -6360 5880 -6300
rect 5940 -6360 6000 -6300
rect 6060 -6360 6120 -6300
rect 6180 -6360 6240 -6300
rect 6300 -6360 6360 -6300
rect 6420 -6360 6480 -6300
rect 6540 -6360 6600 -6300
rect 6660 -6360 6720 -6300
rect 6780 -6360 6840 -6300
rect 6900 -6360 6960 -6300
rect 7020 -6360 7080 -6300
rect 7140 -6360 7200 -6300
rect 7260 -6360 7320 -6300
rect 7380 -6360 7440 -6300
rect 7500 -6360 7560 -6300
rect 7620 -6360 7680 -6300
rect 7740 -6360 7800 -6300
rect 7860 -6360 7920 -6300
rect 7980 -6360 8040 -6300
rect 8100 -6360 8160 -6300
rect 8220 -6360 8280 -6300
rect 8340 -6360 8400 -6300
rect 8460 -6360 8520 -6300
rect 8580 -6360 8640 -6300
rect 8700 -6360 8760 -6300
rect 8820 -6360 8880 -6300
rect 8940 -6360 9000 -6300
rect 9060 -6360 9120 -6300
rect 9180 -6360 9240 -6300
rect 9300 -6360 9360 -6300
rect 9420 -6360 9480 -6300
rect 9540 -6360 9600 -6300
rect 9660 -6360 9720 -6300
rect 9780 -6360 9840 -6300
rect 9900 -6360 9960 -6300
rect 10020 -6360 10080 -6300
rect 10140 -6360 10200 -6300
rect 10260 -6360 10320 -6300
rect 10380 -6360 10440 -6300
rect 10500 -6360 10560 -6300
rect 10620 -6360 10680 -6300
rect 10740 -6360 10800 -6300
rect 10860 -6360 10920 -6300
rect 10980 -6360 11040 -6300
rect 11100 -6360 11160 -6300
rect 11220 -6360 11280 -6300
rect 11340 -6360 11400 -6300
rect 11460 -6360 11520 -6300
rect 11580 -6360 11640 -6300
rect 11700 -6360 11760 -6300
rect 11820 -6360 11880 -6300
rect 11940 -6360 12000 -6300
rect 12060 -6360 12120 -6300
rect 12180 -6360 12240 -6300
rect 12300 -6360 12360 -6300
rect 12420 -6360 12480 -6300
rect 12540 -6360 12600 -6300
rect 12660 -6360 12720 -6300
rect 12780 -6360 12840 -6300
rect 12900 -6360 12960 -6300
rect 13020 -6360 13080 -6300
rect 13140 -6360 13200 -6300
rect 13260 -6360 13320 -6300
rect 13380 -6360 13440 -6300
rect 13500 -6360 13560 -6300
rect 13620 -6360 13680 -6300
rect 13740 -6360 13800 -6300
rect 13860 -6360 13920 -6300
rect 13980 -6360 14040 -6300
rect 14100 -6360 14160 -6300
rect 14220 -6360 14280 -6300
rect 14340 -6360 14400 -6300
rect 14460 -6360 14520 -6300
rect 14580 -6360 14640 -6300
rect 14700 -6360 14760 -6300
rect 14820 -6360 14880 -6300
rect 14940 -6360 15000 -6300
rect 15060 -6360 15120 -6300
rect 15180 -6360 15240 -6300
rect 15300 -6360 15360 -6300
rect 15420 -6360 15480 -6300
rect 15540 -6360 15600 -6300
rect 15660 -6360 15720 -6300
rect 15780 -6360 15840 -6300
rect 15900 -6360 15960 -6300
rect 16020 -6360 16080 -6300
rect 16140 -6360 16200 -6300
rect 16260 -6360 16320 -6300
rect 16380 -6360 16440 -6300
rect 16500 -6360 16560 -6300
rect 16620 -6360 16680 -6300
rect 16740 -6360 16800 -6300
rect 16860 -6360 16920 -6300
rect 16980 -6360 17040 -6300
rect 17100 -6360 17160 -6300
rect 17220 -6360 17280 -6300
rect 17340 -6360 17400 -6300
rect 17460 -6360 17520 -6300
rect 17580 -6360 17640 -6300
rect 17700 -6360 17760 -6300
rect 17820 -6360 17880 -6300
rect 17940 -6360 18000 -6300
rect 18060 -6360 18120 -6300
rect 18180 -6360 18240 -6300
rect 18300 -6360 18360 -6300
rect 18420 -6360 18480 -6300
rect 18540 -6360 18600 -6300
rect 18660 -6360 18720 -6300
rect 18780 -6360 18840 -6300
rect 18900 -6360 18960 -6300
rect 19020 -6360 19080 -6300
rect 19140 -6360 19200 -6300
rect 19260 -6360 19320 -6300
rect 19380 -6360 19440 -6300
rect 19500 -6360 19560 -6300
rect 19620 -6360 19680 -6300
rect 19740 -6360 19800 -6300
rect 19860 -6360 19920 -6300
rect 19980 -6360 20040 -6300
<< locali >>
rect -20 0 60 60
rect 120 0 180 60
rect 240 0 300 60
rect 360 0 420 60
rect 480 0 540 60
rect 600 0 660 60
rect 720 0 780 60
rect 840 0 900 60
rect 960 0 1020 60
rect 1080 0 1140 60
rect 1200 0 1260 60
rect 1320 0 1380 60
rect 1440 0 1500 60
rect 1560 0 1620 60
rect 1680 0 1740 60
rect 1800 0 1860 60
rect 1920 0 1980 60
rect 2040 0 2100 60
rect 2160 0 2220 60
rect 2280 0 2340 60
rect 2400 0 2460 60
rect 2520 0 2580 60
rect 2640 0 2700 60
rect 2760 0 2820 60
rect 2880 0 2940 60
rect 3000 0 3060 60
rect 3120 0 3180 60
rect 3240 0 3300 60
rect 3360 0 3420 60
rect 3480 0 3540 60
rect 3600 0 3660 60
rect 3720 0 3780 60
rect 3840 0 3900 60
rect 3960 0 4020 60
rect 4080 0 4140 60
rect 4200 0 4260 60
rect 4320 0 4380 60
rect 4440 0 4500 60
rect 4560 0 4620 60
rect 4680 0 4740 60
rect 4800 0 4860 60
rect 4920 0 4980 60
rect 5040 0 5100 60
rect 5160 0 5220 60
rect 5280 0 5340 60
rect 5400 0 5460 60
rect 5520 0 5580 60
rect 5640 0 5700 60
rect 5760 0 5820 60
rect 5880 0 5940 60
rect 6000 0 6060 60
rect 6120 0 6180 60
rect 6240 0 6300 60
rect 6360 0 6420 60
rect 6480 0 6540 60
rect 6600 0 6660 60
rect 6720 0 6780 60
rect 6840 0 6900 60
rect 6960 0 7020 60
rect 7080 0 7140 60
rect 7200 0 7260 60
rect 7320 0 7380 60
rect 7440 0 7500 60
rect 7560 0 7620 60
rect 7680 0 7740 60
rect 7800 0 7860 60
rect 7920 0 7980 60
rect 8040 0 8100 60
rect 8160 0 8220 60
rect 8280 0 8340 60
rect 8400 0 8460 60
rect 8520 0 8580 60
rect 8640 0 8700 60
rect 8760 0 8820 60
rect 8880 0 8940 60
rect 9000 0 9060 60
rect 9120 0 9180 60
rect 9240 0 9300 60
rect 9360 0 9420 60
rect 9480 0 9540 60
rect 9600 0 9660 60
rect 9720 0 9780 60
rect 9840 0 9900 60
rect 9960 0 10020 60
rect 10080 0 10140 60
rect 10200 0 10260 60
rect 10320 0 10380 60
rect 10440 0 10500 60
rect 10560 0 10620 60
rect 10680 0 10740 60
rect 10800 0 10860 60
rect 10920 0 10980 60
rect 11040 0 11100 60
rect 11160 0 11220 60
rect 11280 0 11340 60
rect 11400 0 11460 60
rect 11520 0 11580 60
rect 11640 0 11700 60
rect 11760 0 11820 60
rect 11880 0 11940 60
rect 12000 0 12060 60
rect 12120 0 12180 60
rect 12240 0 12300 60
rect 12360 0 12420 60
rect 12480 0 12540 60
rect 12600 0 12660 60
rect 12720 0 12780 60
rect 12840 0 12900 60
rect 12960 0 13020 60
rect 13080 0 13140 60
rect 13200 0 13260 60
rect 13320 0 13380 60
rect 13440 0 13500 60
rect 13560 0 13620 60
rect 13680 0 13740 60
rect 13800 0 13860 60
rect 13920 0 13980 60
rect 14040 0 14100 60
rect 14160 0 14220 60
rect 14280 0 14340 60
rect 14400 0 14460 60
rect 14520 0 14580 60
rect 14640 0 14700 60
rect 14760 0 14820 60
rect 14880 0 14940 60
rect 15000 0 15060 60
rect 15120 0 15180 60
rect 15240 0 15300 60
rect 15360 0 15420 60
rect 15480 0 15540 60
rect 15600 0 15660 60
rect 15720 0 15780 60
rect 15840 0 15900 60
rect 15960 0 16020 60
rect 16080 0 16140 60
rect 16200 0 16260 60
rect 16320 0 16380 60
rect 16440 0 16500 60
rect 16560 0 16620 60
rect 16680 0 16740 60
rect 16800 0 16860 60
rect 16920 0 16980 60
rect 17040 0 17100 60
rect 17160 0 17220 60
rect 17280 0 17340 60
rect 17400 0 17460 60
rect 17520 0 17580 60
rect 17640 0 17700 60
rect 17760 0 17820 60
rect 17880 0 17940 60
rect 18000 0 18060 60
rect -20 -40 40 0
rect -20 -160 40 -100
rect -20 -280 40 -220
rect -20 -400 40 -340
rect -20 -520 40 -460
rect -20 -640 40 -580
rect -20 -760 40 -700
rect -20 -880 40 -820
rect -20 -1000 40 -940
rect -20 -1120 40 -1060
rect -20 -1240 40 -1180
rect -20 -1360 40 -1300
rect -20 -1480 40 -1420
rect -20 -1600 40 -1540
rect -20 -1720 40 -1660
rect -20 -1840 40 -1780
rect -20 -1960 40 -1900
rect -20 -2080 40 -2020
rect -20 -2200 40 -2140
rect -20 -2320 40 -2260
rect -20 -2440 40 -2380
rect -20 -2560 40 -2500
rect -20 -2680 40 -2620
rect -20 -2800 40 -2740
rect -20 -2920 40 -2860
rect -20 -3020 40 -2980
rect -1680 -3186 -1640 -3126
rect -1580 -3186 -1520 -3126
rect -1460 -3186 -1400 -3126
rect -1340 -3186 -1280 -3126
rect -1220 -3186 -1160 -3126
rect -1100 -3186 -1040 -3126
rect -980 -3186 -920 -3126
rect -860 -3186 -800 -3126
rect -740 -3186 -680 -3126
rect -620 -3186 -560 -3126
rect -500 -3186 -440 -3126
rect -380 -3186 -320 -3126
rect -260 -3186 -200 -3126
rect -140 -3186 -80 -3126
rect -20 -3186 40 -3080
rect 18120 -40 18180 60
rect 18120 -160 18180 -100
rect 18120 -280 18180 -220
rect 18120 -400 18180 -340
rect 18120 -520 18180 -460
rect 18120 -640 18180 -580
rect 18120 -760 18180 -700
rect 18120 -880 18180 -820
rect 18120 -1000 18180 -940
rect 18120 -1120 18180 -1060
rect 18120 -1240 18180 -1180
rect 18120 -1360 18180 -1300
rect 18120 -1480 18180 -1420
rect 18120 -1600 18180 -1540
rect 18120 -1720 18180 -1660
rect 18120 -1840 18180 -1780
rect 18120 -1960 18180 -1900
rect 18120 -2080 18180 -2020
rect 18120 -2200 18180 -2140
rect 18120 -2320 18180 -2260
rect 18120 -2440 18180 -2380
rect 18120 -2560 18180 -2500
rect 18120 -2680 18180 -2620
rect 18120 -2800 18180 -2740
rect 18120 -2920 18180 -2860
rect 18120 -3020 18180 -2980
rect 18120 -3126 18180 -3080
rect 100 -3186 140 -3126
rect 200 -3186 260 -3126
rect 320 -3186 380 -3126
rect 440 -3186 500 -3126
rect 560 -3186 620 -3126
rect 680 -3186 740 -3126
rect 800 -3186 860 -3126
rect 920 -3186 980 -3126
rect 1040 -3186 1100 -3126
rect 1160 -3186 1220 -3126
rect 1280 -3186 1340 -3126
rect 1400 -3186 1460 -3126
rect 1520 -3186 1580 -3126
rect 1640 -3186 1700 -3126
rect 1760 -3186 1820 -3126
rect 1880 -3186 1940 -3126
rect 2000 -3186 2060 -3126
rect 2120 -3186 2180 -3126
rect 2240 -3186 2300 -3126
rect 2360 -3186 2420 -3126
rect 2480 -3186 2540 -3126
rect 2600 -3186 2660 -3126
rect 2720 -3186 2780 -3126
rect 2840 -3186 2900 -3126
rect 2960 -3186 3020 -3126
rect 3080 -3186 3140 -3126
rect 3200 -3186 3260 -3126
rect 3320 -3186 3380 -3126
rect 3440 -3186 3500 -3126
rect 3560 -3186 3620 -3126
rect 3680 -3186 3740 -3126
rect 3800 -3186 3860 -3126
rect 3920 -3186 3980 -3126
rect 4040 -3186 4100 -3126
rect 4160 -3186 4220 -3126
rect 4280 -3186 4340 -3126
rect 4400 -3186 4460 -3126
rect 4520 -3186 4580 -3126
rect 4640 -3186 4700 -3126
rect 4760 -3186 4820 -3126
rect 4880 -3186 4940 -3126
rect 5000 -3186 5060 -3126
rect 5120 -3186 5180 -3126
rect 5240 -3186 5300 -3126
rect 5360 -3186 5420 -3126
rect 5480 -3186 5540 -3126
rect 5600 -3186 5660 -3126
rect 5720 -3186 5780 -3126
rect 5840 -3186 5900 -3126
rect 5960 -3186 6020 -3126
rect 6080 -3186 6140 -3126
rect 6200 -3186 6260 -3126
rect 6320 -3186 6380 -3126
rect 6440 -3186 6500 -3126
rect 6560 -3186 6620 -3126
rect 6680 -3186 6740 -3126
rect 6800 -3186 6860 -3126
rect 6920 -3186 6980 -3126
rect 7040 -3186 7100 -3126
rect 7160 -3186 7220 -3126
rect 7280 -3186 7340 -3126
rect 7400 -3186 7460 -3126
rect 7520 -3186 7580 -3126
rect 7640 -3186 7700 -3126
rect 7760 -3186 7820 -3126
rect 7880 -3186 7940 -3126
rect 8000 -3186 8060 -3126
rect 8120 -3186 8180 -3126
rect 8240 -3186 8300 -3126
rect 8360 -3186 8420 -3126
rect 8480 -3186 8540 -3126
rect 8600 -3186 8660 -3126
rect 8720 -3186 8780 -3126
rect 8840 -3186 8900 -3126
rect 8960 -3186 9020 -3126
rect 9080 -3186 9140 -3126
rect 9200 -3186 9260 -3126
rect 9320 -3186 9380 -3126
rect 9440 -3186 9500 -3126
rect 9560 -3186 9620 -3126
rect 9680 -3186 9740 -3126
rect 9800 -3186 9860 -3126
rect 9920 -3186 9980 -3126
rect 10040 -3186 10100 -3126
rect 10160 -3186 10220 -3126
rect 10280 -3186 10340 -3126
rect 10400 -3186 10460 -3126
rect 10520 -3186 10580 -3126
rect 10640 -3186 10700 -3126
rect 10760 -3186 10820 -3126
rect 10880 -3186 10940 -3126
rect 11000 -3186 11060 -3126
rect 11120 -3186 11180 -3126
rect 11240 -3186 11300 -3126
rect 11360 -3186 11420 -3126
rect 11480 -3186 11540 -3126
rect 11600 -3186 11660 -3126
rect 11720 -3186 11780 -3126
rect 11840 -3186 11900 -3126
rect 11960 -3186 12020 -3126
rect 12080 -3186 12140 -3126
rect 12200 -3186 12260 -3126
rect 12320 -3186 12380 -3126
rect 12440 -3186 12500 -3126
rect 12560 -3186 12620 -3126
rect 12680 -3186 12740 -3126
rect 12800 -3186 12860 -3126
rect 12920 -3186 12980 -3126
rect 13040 -3186 13100 -3126
rect 13160 -3186 13220 -3126
rect 13280 -3186 13340 -3126
rect 13400 -3186 13460 -3126
rect 13520 -3186 13580 -3126
rect 13640 -3186 13700 -3126
rect 13760 -3186 13820 -3126
rect 13880 -3186 13940 -3126
rect 14000 -3186 14060 -3126
rect 14120 -3186 14180 -3126
rect 14240 -3186 14300 -3126
rect 14360 -3186 14420 -3126
rect 14480 -3186 14540 -3126
rect 14600 -3186 14660 -3126
rect 14720 -3186 14780 -3126
rect 14840 -3186 14900 -3126
rect 14960 -3186 15020 -3126
rect 15080 -3186 15140 -3126
rect 15200 -3186 15260 -3126
rect 15320 -3186 15380 -3126
rect 15440 -3186 15500 -3126
rect 15560 -3186 15620 -3126
rect 15680 -3186 15740 -3126
rect 15800 -3186 15860 -3126
rect 15920 -3186 15980 -3126
rect 16040 -3186 16100 -3126
rect 16160 -3186 16220 -3126
rect 16280 -3186 16340 -3126
rect 16400 -3186 16460 -3126
rect 16520 -3186 16580 -3126
rect 16640 -3186 16700 -3126
rect 16760 -3186 16820 -3126
rect 16880 -3186 16940 -3126
rect 17000 -3186 17060 -3126
rect 17120 -3186 17180 -3126
rect 17240 -3186 17300 -3126
rect 17360 -3186 17420 -3126
rect 17480 -3186 17540 -3126
rect 17600 -3186 17660 -3126
rect 17720 -3186 17780 -3126
rect 17840 -3186 17900 -3126
rect 17960 -3186 18020 -3126
rect 18080 -3186 18140 -3126
rect 18200 -3186 18260 -3126
rect 18320 -3186 18380 -3126
rect 18440 -3186 18500 -3126
rect 18560 -3186 18620 -3126
rect 18680 -3186 18740 -3126
rect 18800 -3186 18860 -3126
rect 18920 -3186 18980 -3126
rect 19040 -3186 19100 -3126
rect 19160 -3186 19220 -3126
rect 19280 -3186 19340 -3126
rect 19400 -3186 19460 -3126
rect 19520 -3186 19580 -3126
rect 19640 -3186 19700 -3126
rect 19760 -3186 19820 -3126
rect 19880 -3186 19940 -3126
rect 20000 -3186 20060 -3126
rect 20120 -3186 20145 -3126
rect -1680 -3226 -1620 -3186
rect -1680 -3346 -1620 -3286
rect -1680 -3466 -1620 -3406
rect -1680 -3586 -1620 -3526
rect -1680 -3706 -1620 -3646
rect -1680 -3826 -1620 -3766
rect -1680 -3946 -1620 -3886
rect -1680 -4066 -1620 -4006
rect -1680 -4186 -1620 -4126
rect -1680 -4306 -1620 -4246
rect -1680 -4426 -1620 -4366
rect -1680 -4546 -1620 -4486
rect -1680 -4666 -1620 -4606
rect -1680 -4786 -1620 -4726
rect -1680 -4906 -1620 -4846
rect -1680 -5026 -1620 -4966
rect -1680 -5146 -1620 -5086
rect -1680 -5266 -1620 -5206
rect -1680 -5386 -1620 -5326
rect -1680 -5506 -1620 -5446
rect -1680 -5626 -1620 -5566
rect -1680 -5746 -1620 -5686
rect -1680 -5866 -1620 -5806
rect -1680 -5986 -1620 -5926
rect -1680 -6106 -1620 -6046
rect -1680 -6206 -1620 -6166
rect -1680 -6360 -1620 -6266
rect 20080 -3200 20145 -3186
rect 20080 -3246 20140 -3200
rect 20080 -3366 20140 -3306
rect 20080 -3486 20140 -3426
rect 20080 -3606 20140 -3546
rect 20080 -3726 20140 -3666
rect 20080 -3846 20140 -3786
rect 20080 -3966 20140 -3906
rect 20080 -4086 20140 -4026
rect 20080 -4206 20140 -4146
rect 20080 -4326 20140 -4266
rect 20080 -4446 20140 -4386
rect 20080 -4566 20140 -4506
rect 20080 -4686 20140 -4626
rect 20080 -4806 20140 -4746
rect 20080 -4926 20140 -4866
rect 20080 -5046 20140 -4986
rect 20080 -5166 20140 -5106
rect 20080 -5286 20140 -5226
rect 20080 -5406 20140 -5346
rect 20080 -5526 20140 -5466
rect 20080 -5646 20140 -5586
rect 20080 -5766 20140 -5706
rect 20080 -5886 20140 -5826
rect 20080 -6006 20140 -5946
rect 20080 -6126 20140 -6066
rect 20080 -6240 20140 -6186
rect -1560 -6360 -1500 -6300
rect -1440 -6360 -1380 -6300
rect -1320 -6360 -1260 -6300
rect -1200 -6360 -1140 -6300
rect -1080 -6360 -1020 -6300
rect -960 -6360 -900 -6300
rect -840 -6360 -780 -6300
rect -720 -6360 -660 -6300
rect -600 -6360 -540 -6300
rect -480 -6360 -420 -6300
rect -360 -6360 -300 -6300
rect -240 -6360 -180 -6300
rect -120 -6360 -60 -6300
rect 0 -6360 60 -6300
rect 120 -6360 180 -6300
rect 240 -6360 300 -6300
rect 360 -6360 420 -6300
rect 480 -6360 540 -6300
rect 600 -6360 660 -6300
rect 720 -6360 780 -6300
rect 840 -6360 900 -6300
rect 960 -6360 1020 -6300
rect 1080 -6360 1140 -6300
rect 1200 -6360 1260 -6300
rect 1320 -6360 1380 -6300
rect 1440 -6360 1500 -6300
rect 1560 -6360 1620 -6300
rect 1680 -6360 1740 -6300
rect 1800 -6360 1860 -6300
rect 1920 -6360 1980 -6300
rect 2040 -6360 2100 -6300
rect 2160 -6360 2220 -6300
rect 2280 -6360 2340 -6300
rect 2400 -6360 2460 -6300
rect 2520 -6360 2580 -6300
rect 2640 -6360 2700 -6300
rect 2760 -6360 2820 -6300
rect 2880 -6360 2940 -6300
rect 3000 -6360 3060 -6300
rect 3120 -6360 3180 -6300
rect 3240 -6360 3300 -6300
rect 3360 -6360 3420 -6300
rect 3480 -6360 3540 -6300
rect 3600 -6360 3660 -6300
rect 3720 -6360 3780 -6300
rect 3840 -6360 3900 -6300
rect 3960 -6360 4020 -6300
rect 4080 -6360 4140 -6300
rect 4200 -6360 4260 -6300
rect 4320 -6360 4380 -6300
rect 4440 -6360 4500 -6300
rect 4560 -6360 4620 -6300
rect 4680 -6360 4740 -6300
rect 4800 -6360 4860 -6300
rect 4920 -6360 4980 -6300
rect 5040 -6360 5100 -6300
rect 5160 -6360 5220 -6300
rect 5280 -6360 5340 -6300
rect 5400 -6360 5460 -6300
rect 5520 -6360 5580 -6300
rect 5640 -6360 5700 -6300
rect 5760 -6360 5820 -6300
rect 5880 -6360 5940 -6300
rect 6000 -6360 6060 -6300
rect 6120 -6360 6180 -6300
rect 6240 -6360 6300 -6300
rect 6360 -6360 6420 -6300
rect 6480 -6360 6540 -6300
rect 6600 -6360 6660 -6300
rect 6720 -6360 6780 -6300
rect 6840 -6360 6900 -6300
rect 6960 -6360 7020 -6300
rect 7080 -6360 7140 -6300
rect 7200 -6360 7260 -6300
rect 7320 -6360 7380 -6300
rect 7440 -6360 7500 -6300
rect 7560 -6360 7620 -6300
rect 7680 -6360 7740 -6300
rect 7800 -6360 7860 -6300
rect 7920 -6360 7980 -6300
rect 8040 -6360 8100 -6300
rect 8160 -6360 8220 -6300
rect 8280 -6360 8340 -6300
rect 8400 -6360 8460 -6300
rect 8520 -6360 8580 -6300
rect 8640 -6360 8700 -6300
rect 8760 -6360 8820 -6300
rect 8880 -6360 8940 -6300
rect 9000 -6360 9060 -6300
rect 9120 -6360 9180 -6300
rect 9240 -6360 9300 -6300
rect 9360 -6360 9420 -6300
rect 9480 -6360 9540 -6300
rect 9600 -6360 9660 -6300
rect 9720 -6360 9780 -6300
rect 9840 -6360 9900 -6300
rect 9960 -6360 10020 -6300
rect 10080 -6360 10140 -6300
rect 10200 -6360 10260 -6300
rect 10320 -6360 10380 -6300
rect 10440 -6360 10500 -6300
rect 10560 -6360 10620 -6300
rect 10680 -6360 10740 -6300
rect 10800 -6360 10860 -6300
rect 10920 -6360 10980 -6300
rect 11040 -6360 11100 -6300
rect 11160 -6360 11220 -6300
rect 11280 -6360 11340 -6300
rect 11400 -6360 11460 -6300
rect 11520 -6360 11580 -6300
rect 11640 -6360 11700 -6300
rect 11760 -6360 11820 -6300
rect 11880 -6360 11940 -6300
rect 12000 -6360 12060 -6300
rect 12120 -6360 12180 -6300
rect 12240 -6360 12300 -6300
rect 12360 -6360 12420 -6300
rect 12480 -6360 12540 -6300
rect 12600 -6360 12660 -6300
rect 12720 -6360 12780 -6300
rect 12840 -6360 12900 -6300
rect 12960 -6360 13020 -6300
rect 13080 -6360 13140 -6300
rect 13200 -6360 13260 -6300
rect 13320 -6360 13380 -6300
rect 13440 -6360 13500 -6300
rect 13560 -6360 13620 -6300
rect 13680 -6360 13740 -6300
rect 13800 -6360 13860 -6300
rect 13920 -6360 13980 -6300
rect 14040 -6360 14100 -6300
rect 14160 -6360 14220 -6300
rect 14280 -6360 14340 -6300
rect 14400 -6360 14460 -6300
rect 14520 -6360 14580 -6300
rect 14640 -6360 14700 -6300
rect 14760 -6360 14820 -6300
rect 14880 -6360 14940 -6300
rect 15000 -6360 15060 -6300
rect 15120 -6360 15180 -6300
rect 15240 -6360 15300 -6300
rect 15360 -6360 15420 -6300
rect 15480 -6360 15540 -6300
rect 15600 -6360 15660 -6300
rect 15720 -6360 15780 -6300
rect 15840 -6360 15900 -6300
rect 15960 -6360 16020 -6300
rect 16080 -6360 16140 -6300
rect 16200 -6360 16260 -6300
rect 16320 -6360 16380 -6300
rect 16440 -6360 16500 -6300
rect 16560 -6360 16620 -6300
rect 16680 -6360 16740 -6300
rect 16800 -6360 16860 -6300
rect 16920 -6360 16980 -6300
rect 17040 -6360 17100 -6300
rect 17160 -6360 17220 -6300
rect 17280 -6360 17340 -6300
rect 17400 -6360 17460 -6300
rect 17520 -6360 17580 -6300
rect 17640 -6360 17700 -6300
rect 17760 -6360 17820 -6300
rect 17880 -6360 17940 -6300
rect 18000 -6360 18060 -6300
rect 18120 -6360 18180 -6300
rect 18240 -6360 18300 -6300
rect 18360 -6360 18420 -6300
rect 18480 -6360 18540 -6300
rect 18600 -6360 18660 -6300
rect 18720 -6360 18780 -6300
rect 18840 -6360 18900 -6300
rect 18960 -6360 19020 -6300
rect 19080 -6360 19140 -6300
rect 19200 -6360 19260 -6300
rect 19320 -6360 19380 -6300
rect 19440 -6360 19500 -6300
rect 19560 -6360 19620 -6300
rect 19680 -6360 19740 -6300
rect 19800 -6360 19860 -6300
rect 19920 -6360 19980 -6300
rect 20040 -6360 20140 -6300
<< end >>
