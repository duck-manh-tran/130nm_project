magic
tech sky130A
timestamp 1623530672
<< metal3 >>
rect 0 10480 12200 10500
rect 0 10440 20 10480
rect 60 10440 80 10480
rect 120 10440 140 10480
rect 180 10440 1820 10480
rect 1860 10440 1880 10480
rect 1920 10440 1940 10480
rect 1980 10440 4620 10480
rect 4660 10440 4680 10480
rect 4720 10440 4740 10480
rect 4780 10440 7420 10480
rect 7460 10440 7480 10480
rect 7520 10440 7540 10480
rect 7580 10440 10220 10480
rect 10260 10440 10280 10480
rect 10320 10440 10340 10480
rect 10380 10440 12020 10480
rect 12060 10440 12080 10480
rect 12120 10440 12140 10480
rect 12180 10440 12200 10480
rect 0 10420 12200 10440
rect 0 10380 20 10420
rect 60 10380 80 10420
rect 120 10380 140 10420
rect 180 10380 1820 10420
rect 1860 10380 1880 10420
rect 1920 10380 1940 10420
rect 1980 10380 4620 10420
rect 4660 10380 4680 10420
rect 4720 10380 4740 10420
rect 4780 10380 7420 10420
rect 7460 10380 7480 10420
rect 7520 10380 7540 10420
rect 7580 10380 10220 10420
rect 10260 10380 10280 10420
rect 10320 10380 10340 10420
rect 10380 10380 12020 10420
rect 12060 10380 12080 10420
rect 12120 10380 12140 10420
rect 12180 10380 12200 10420
rect 0 10360 12200 10380
rect 0 10320 20 10360
rect 60 10320 80 10360
rect 120 10320 140 10360
rect 180 10320 1820 10360
rect 1860 10320 1880 10360
rect 1920 10320 1940 10360
rect 1980 10320 4620 10360
rect 4660 10320 4680 10360
rect 4720 10320 4740 10360
rect 4780 10320 7420 10360
rect 7460 10320 7480 10360
rect 7520 10320 7540 10360
rect 7580 10320 10220 10360
rect 10260 10320 10280 10360
rect 10320 10320 10340 10360
rect 10380 10320 12020 10360
rect 12060 10320 12080 10360
rect 12120 10320 12140 10360
rect 12180 10320 12200 10360
rect 0 10300 12200 10320
rect 400 10080 11800 10100
rect 400 10040 420 10080
rect 460 10040 480 10080
rect 520 10040 540 10080
rect 580 10040 3220 10080
rect 3260 10040 3280 10080
rect 3320 10040 3340 10080
rect 3380 10040 6020 10080
rect 6060 10040 6080 10080
rect 6120 10040 6140 10080
rect 6180 10040 8820 10080
rect 8860 10040 8880 10080
rect 8920 10040 8940 10080
rect 8980 10040 11620 10080
rect 11660 10040 11680 10080
rect 11720 10040 11740 10080
rect 11780 10040 11800 10080
rect 400 10020 11800 10040
rect 400 9980 420 10020
rect 460 9980 480 10020
rect 520 9980 540 10020
rect 580 9980 3220 10020
rect 3260 9980 3280 10020
rect 3320 9980 3340 10020
rect 3380 9980 6020 10020
rect 6060 9980 6080 10020
rect 6120 9980 6140 10020
rect 6180 9980 8820 10020
rect 8860 9980 8880 10020
rect 8920 9980 8940 10020
rect 8980 9980 11620 10020
rect 11660 9980 11680 10020
rect 11720 9980 11740 10020
rect 11780 9980 11800 10020
rect 400 9960 11800 9980
rect 400 9920 420 9960
rect 460 9920 480 9960
rect 520 9920 540 9960
rect 580 9920 3220 9960
rect 3260 9920 3280 9960
rect 3320 9920 3340 9960
rect 3380 9920 6020 9960
rect 6060 9920 6080 9960
rect 6120 9920 6140 9960
rect 6180 9920 8820 9960
rect 8860 9920 8880 9960
rect 8920 9920 8940 9960
rect 8980 9920 11620 9960
rect 11660 9920 11680 9960
rect 11720 9920 11740 9960
rect 11780 9920 11800 9960
rect 400 9900 11800 9920
rect 400 580 11800 600
rect 400 540 420 580
rect 460 540 480 580
rect 520 540 540 580
rect 580 540 3220 580
rect 3260 540 3280 580
rect 3320 540 3340 580
rect 3380 540 6020 580
rect 6060 540 6080 580
rect 6120 540 6140 580
rect 6180 540 8820 580
rect 8860 540 8880 580
rect 8920 540 8940 580
rect 8980 540 11620 580
rect 11660 540 11680 580
rect 11720 540 11740 580
rect 11780 540 11800 580
rect 400 520 11800 540
rect 400 480 420 520
rect 460 480 480 520
rect 520 480 540 520
rect 580 480 3220 520
rect 3260 480 3280 520
rect 3320 480 3340 520
rect 3380 480 6020 520
rect 6060 480 6080 520
rect 6120 480 6140 520
rect 6180 480 8820 520
rect 8860 480 8880 520
rect 8920 480 8940 520
rect 8980 480 11620 520
rect 11660 480 11680 520
rect 11720 480 11740 520
rect 11780 480 11800 520
rect 400 460 11800 480
rect 400 420 420 460
rect 460 420 480 460
rect 520 420 540 460
rect 580 420 3220 460
rect 3260 420 3280 460
rect 3320 420 3340 460
rect 3380 420 6020 460
rect 6060 420 6080 460
rect 6120 420 6140 460
rect 6180 420 8820 460
rect 8860 420 8880 460
rect 8920 420 8940 460
rect 8980 420 11620 460
rect 11660 420 11680 460
rect 11720 420 11740 460
rect 11780 420 11800 460
rect 400 400 11800 420
rect 0 180 12200 200
rect 0 140 20 180
rect 60 140 80 180
rect 120 140 140 180
rect 180 140 1820 180
rect 1860 140 1880 180
rect 1920 140 1940 180
rect 1980 140 4620 180
rect 4660 140 4680 180
rect 4720 140 4740 180
rect 4780 140 7420 180
rect 7460 140 7480 180
rect 7520 140 7540 180
rect 7580 140 10220 180
rect 10260 140 10280 180
rect 10320 140 10340 180
rect 10380 140 12020 180
rect 12060 140 12080 180
rect 12120 140 12140 180
rect 12180 140 12200 180
rect 0 120 12200 140
rect 0 80 20 120
rect 60 80 80 120
rect 120 80 140 120
rect 180 80 1820 120
rect 1860 80 1880 120
rect 1920 80 1940 120
rect 1980 80 4620 120
rect 4660 80 4680 120
rect 4720 80 4740 120
rect 4780 80 7420 120
rect 7460 80 7480 120
rect 7520 80 7540 120
rect 7580 80 10220 120
rect 10260 80 10280 120
rect 10320 80 10340 120
rect 10380 80 12020 120
rect 12060 80 12080 120
rect 12120 80 12140 120
rect 12180 80 12200 120
rect 0 60 12200 80
rect 0 20 20 60
rect 60 20 80 60
rect 120 20 140 60
rect 180 20 1820 60
rect 1860 20 1880 60
rect 1920 20 1940 60
rect 1980 20 4620 60
rect 4660 20 4680 60
rect 4720 20 4740 60
rect 4780 20 7420 60
rect 7460 20 7480 60
rect 7520 20 7540 60
rect 7580 20 10220 60
rect 10260 20 10280 60
rect 10320 20 10340 60
rect 10380 20 12020 60
rect 12060 20 12080 60
rect 12120 20 12140 60
rect 12180 20 12200 60
rect 0 0 12200 20
<< via3 >>
rect 20 10440 60 10480
rect 80 10440 120 10480
rect 140 10440 180 10480
rect 1820 10440 1860 10480
rect 1880 10440 1920 10480
rect 1940 10440 1980 10480
rect 4620 10440 4660 10480
rect 4680 10440 4720 10480
rect 4740 10440 4780 10480
rect 7420 10440 7460 10480
rect 7480 10440 7520 10480
rect 7540 10440 7580 10480
rect 10220 10440 10260 10480
rect 10280 10440 10320 10480
rect 10340 10440 10380 10480
rect 12020 10440 12060 10480
rect 12080 10440 12120 10480
rect 12140 10440 12180 10480
rect 20 10380 60 10420
rect 80 10380 120 10420
rect 140 10380 180 10420
rect 1820 10380 1860 10420
rect 1880 10380 1920 10420
rect 1940 10380 1980 10420
rect 4620 10380 4660 10420
rect 4680 10380 4720 10420
rect 4740 10380 4780 10420
rect 7420 10380 7460 10420
rect 7480 10380 7520 10420
rect 7540 10380 7580 10420
rect 10220 10380 10260 10420
rect 10280 10380 10320 10420
rect 10340 10380 10380 10420
rect 12020 10380 12060 10420
rect 12080 10380 12120 10420
rect 12140 10380 12180 10420
rect 20 10320 60 10360
rect 80 10320 120 10360
rect 140 10320 180 10360
rect 1820 10320 1860 10360
rect 1880 10320 1920 10360
rect 1940 10320 1980 10360
rect 4620 10320 4660 10360
rect 4680 10320 4720 10360
rect 4740 10320 4780 10360
rect 7420 10320 7460 10360
rect 7480 10320 7520 10360
rect 7540 10320 7580 10360
rect 10220 10320 10260 10360
rect 10280 10320 10320 10360
rect 10340 10320 10380 10360
rect 12020 10320 12060 10360
rect 12080 10320 12120 10360
rect 12140 10320 12180 10360
rect 420 10040 460 10080
rect 480 10040 520 10080
rect 540 10040 580 10080
rect 3220 10040 3260 10080
rect 3280 10040 3320 10080
rect 3340 10040 3380 10080
rect 6020 10040 6060 10080
rect 6080 10040 6120 10080
rect 6140 10040 6180 10080
rect 8820 10040 8860 10080
rect 8880 10040 8920 10080
rect 8940 10040 8980 10080
rect 11620 10040 11660 10080
rect 11680 10040 11720 10080
rect 11740 10040 11780 10080
rect 420 9980 460 10020
rect 480 9980 520 10020
rect 540 9980 580 10020
rect 3220 9980 3260 10020
rect 3280 9980 3320 10020
rect 3340 9980 3380 10020
rect 6020 9980 6060 10020
rect 6080 9980 6120 10020
rect 6140 9980 6180 10020
rect 8820 9980 8860 10020
rect 8880 9980 8920 10020
rect 8940 9980 8980 10020
rect 11620 9980 11660 10020
rect 11680 9980 11720 10020
rect 11740 9980 11780 10020
rect 420 9920 460 9960
rect 480 9920 520 9960
rect 540 9920 580 9960
rect 3220 9920 3260 9960
rect 3280 9920 3320 9960
rect 3340 9920 3380 9960
rect 6020 9920 6060 9960
rect 6080 9920 6120 9960
rect 6140 9920 6180 9960
rect 8820 9920 8860 9960
rect 8880 9920 8920 9960
rect 8940 9920 8980 9960
rect 11620 9920 11660 9960
rect 11680 9920 11720 9960
rect 11740 9920 11780 9960
rect 420 540 460 580
rect 480 540 520 580
rect 540 540 580 580
rect 3220 540 3260 580
rect 3280 540 3320 580
rect 3340 540 3380 580
rect 6020 540 6060 580
rect 6080 540 6120 580
rect 6140 540 6180 580
rect 8820 540 8860 580
rect 8880 540 8920 580
rect 8940 540 8980 580
rect 11620 540 11660 580
rect 11680 540 11720 580
rect 11740 540 11780 580
rect 420 480 460 520
rect 480 480 520 520
rect 540 480 580 520
rect 3220 480 3260 520
rect 3280 480 3320 520
rect 3340 480 3380 520
rect 6020 480 6060 520
rect 6080 480 6120 520
rect 6140 480 6180 520
rect 8820 480 8860 520
rect 8880 480 8920 520
rect 8940 480 8980 520
rect 11620 480 11660 520
rect 11680 480 11720 520
rect 11740 480 11780 520
rect 420 420 460 460
rect 480 420 520 460
rect 540 420 580 460
rect 3220 420 3260 460
rect 3280 420 3320 460
rect 3340 420 3380 460
rect 6020 420 6060 460
rect 6080 420 6120 460
rect 6140 420 6180 460
rect 8820 420 8860 460
rect 8880 420 8920 460
rect 8940 420 8980 460
rect 11620 420 11660 460
rect 11680 420 11720 460
rect 11740 420 11780 460
rect 20 140 60 180
rect 80 140 120 180
rect 140 140 180 180
rect 1820 140 1860 180
rect 1880 140 1920 180
rect 1940 140 1980 180
rect 4620 140 4660 180
rect 4680 140 4720 180
rect 4740 140 4780 180
rect 7420 140 7460 180
rect 7480 140 7520 180
rect 7540 140 7580 180
rect 10220 140 10260 180
rect 10280 140 10320 180
rect 10340 140 10380 180
rect 12020 140 12060 180
rect 12080 140 12120 180
rect 12140 140 12180 180
rect 20 80 60 120
rect 80 80 120 120
rect 140 80 180 120
rect 1820 80 1860 120
rect 1880 80 1920 120
rect 1940 80 1980 120
rect 4620 80 4660 120
rect 4680 80 4720 120
rect 4740 80 4780 120
rect 7420 80 7460 120
rect 7480 80 7520 120
rect 7540 80 7580 120
rect 10220 80 10260 120
rect 10280 80 10320 120
rect 10340 80 10380 120
rect 12020 80 12060 120
rect 12080 80 12120 120
rect 12140 80 12180 120
rect 20 20 60 60
rect 80 20 120 60
rect 140 20 180 60
rect 1820 20 1860 60
rect 1880 20 1920 60
rect 1940 20 1980 60
rect 4620 20 4660 60
rect 4680 20 4720 60
rect 4740 20 4780 60
rect 7420 20 7460 60
rect 7480 20 7520 60
rect 7540 20 7580 60
rect 10220 20 10260 60
rect 10280 20 10320 60
rect 10340 20 10380 60
rect 12020 20 12060 60
rect 12080 20 12120 60
rect 12140 20 12180 60
<< metal4 >>
rect 0 10480 200 10500
rect 0 10440 20 10480
rect 60 10440 80 10480
rect 120 10440 140 10480
rect 180 10440 200 10480
rect 0 10420 200 10440
rect 0 10380 20 10420
rect 60 10380 80 10420
rect 120 10380 140 10420
rect 180 10380 200 10420
rect 0 10360 200 10380
rect 0 10320 20 10360
rect 60 10320 80 10360
rect 120 10320 140 10360
rect 180 10320 200 10360
rect 0 180 200 10320
rect 1800 10480 2000 10500
rect 1800 10440 1820 10480
rect 1860 10440 1880 10480
rect 1920 10440 1940 10480
rect 1980 10440 2000 10480
rect 1800 10420 2000 10440
rect 1800 10380 1820 10420
rect 1860 10380 1880 10420
rect 1920 10380 1940 10420
rect 1980 10380 2000 10420
rect 1800 10360 2000 10380
rect 1800 10320 1820 10360
rect 1860 10320 1880 10360
rect 1920 10320 1940 10360
rect 1980 10320 2000 10360
rect 400 10080 600 10100
rect 400 10040 420 10080
rect 460 10040 480 10080
rect 520 10040 540 10080
rect 580 10040 600 10080
rect 400 10020 600 10040
rect 400 9980 420 10020
rect 460 9980 480 10020
rect 520 9980 540 10020
rect 580 9980 600 10020
rect 400 9960 600 9980
rect 400 9920 420 9960
rect 460 9920 480 9960
rect 520 9920 540 9960
rect 580 9920 600 9960
rect 400 580 600 9920
rect 400 540 420 580
rect 460 540 480 580
rect 520 540 540 580
rect 580 540 600 580
rect 400 520 600 540
rect 400 480 420 520
rect 460 480 480 520
rect 520 480 540 520
rect 580 480 600 520
rect 400 460 600 480
rect 400 420 420 460
rect 460 420 480 460
rect 520 420 540 460
rect 580 420 600 460
rect 400 400 600 420
rect 0 140 20 180
rect 60 140 80 180
rect 120 140 140 180
rect 180 140 200 180
rect 0 120 200 140
rect 0 80 20 120
rect 60 80 80 120
rect 120 80 140 120
rect 180 80 200 120
rect 0 60 200 80
rect 0 20 20 60
rect 60 20 80 60
rect 120 20 140 60
rect 180 20 200 60
rect 0 0 200 20
rect 1800 180 2000 10320
rect 4600 10480 4800 10500
rect 4600 10440 4620 10480
rect 4660 10440 4680 10480
rect 4720 10440 4740 10480
rect 4780 10440 4800 10480
rect 4600 10420 4800 10440
rect 4600 10380 4620 10420
rect 4660 10380 4680 10420
rect 4720 10380 4740 10420
rect 4780 10380 4800 10420
rect 4600 10360 4800 10380
rect 4600 10320 4620 10360
rect 4660 10320 4680 10360
rect 4720 10320 4740 10360
rect 4780 10320 4800 10360
rect 3200 10080 3400 10100
rect 3200 10040 3220 10080
rect 3260 10040 3280 10080
rect 3320 10040 3340 10080
rect 3380 10040 3400 10080
rect 3200 10020 3400 10040
rect 3200 9980 3220 10020
rect 3260 9980 3280 10020
rect 3320 9980 3340 10020
rect 3380 9980 3400 10020
rect 3200 9960 3400 9980
rect 3200 9920 3220 9960
rect 3260 9920 3280 9960
rect 3320 9920 3340 9960
rect 3380 9920 3400 9960
rect 3200 580 3400 9920
rect 3200 540 3220 580
rect 3260 540 3280 580
rect 3320 540 3340 580
rect 3380 540 3400 580
rect 3200 520 3400 540
rect 3200 480 3220 520
rect 3260 480 3280 520
rect 3320 480 3340 520
rect 3380 480 3400 520
rect 3200 460 3400 480
rect 3200 420 3220 460
rect 3260 420 3280 460
rect 3320 420 3340 460
rect 3380 420 3400 460
rect 3200 400 3400 420
rect 1800 140 1820 180
rect 1860 140 1880 180
rect 1920 140 1940 180
rect 1980 140 2000 180
rect 1800 120 2000 140
rect 1800 80 1820 120
rect 1860 80 1880 120
rect 1920 80 1940 120
rect 1980 80 2000 120
rect 1800 60 2000 80
rect 1800 20 1820 60
rect 1860 20 1880 60
rect 1920 20 1940 60
rect 1980 20 2000 60
rect 1800 0 2000 20
rect 4600 180 4800 10320
rect 7400 10480 7600 10500
rect 7400 10440 7420 10480
rect 7460 10440 7480 10480
rect 7520 10440 7540 10480
rect 7580 10440 7600 10480
rect 7400 10420 7600 10440
rect 7400 10380 7420 10420
rect 7460 10380 7480 10420
rect 7520 10380 7540 10420
rect 7580 10380 7600 10420
rect 7400 10360 7600 10380
rect 7400 10320 7420 10360
rect 7460 10320 7480 10360
rect 7520 10320 7540 10360
rect 7580 10320 7600 10360
rect 6000 10080 6200 10100
rect 6000 10040 6020 10080
rect 6060 10040 6080 10080
rect 6120 10040 6140 10080
rect 6180 10040 6200 10080
rect 6000 10020 6200 10040
rect 6000 9980 6020 10020
rect 6060 9980 6080 10020
rect 6120 9980 6140 10020
rect 6180 9980 6200 10020
rect 6000 9960 6200 9980
rect 6000 9920 6020 9960
rect 6060 9920 6080 9960
rect 6120 9920 6140 9960
rect 6180 9920 6200 9960
rect 6000 580 6200 9920
rect 6000 540 6020 580
rect 6060 540 6080 580
rect 6120 540 6140 580
rect 6180 540 6200 580
rect 6000 520 6200 540
rect 6000 480 6020 520
rect 6060 480 6080 520
rect 6120 480 6140 520
rect 6180 480 6200 520
rect 6000 460 6200 480
rect 6000 420 6020 460
rect 6060 420 6080 460
rect 6120 420 6140 460
rect 6180 420 6200 460
rect 6000 400 6200 420
rect 4600 140 4620 180
rect 4660 140 4680 180
rect 4720 140 4740 180
rect 4780 140 4800 180
rect 4600 120 4800 140
rect 4600 80 4620 120
rect 4660 80 4680 120
rect 4720 80 4740 120
rect 4780 80 4800 120
rect 4600 60 4800 80
rect 4600 20 4620 60
rect 4660 20 4680 60
rect 4720 20 4740 60
rect 4780 20 4800 60
rect 4600 0 4800 20
rect 7400 180 7600 10320
rect 10200 10480 10400 10500
rect 10200 10440 10220 10480
rect 10260 10440 10280 10480
rect 10320 10440 10340 10480
rect 10380 10440 10400 10480
rect 10200 10420 10400 10440
rect 10200 10380 10220 10420
rect 10260 10380 10280 10420
rect 10320 10380 10340 10420
rect 10380 10380 10400 10420
rect 10200 10360 10400 10380
rect 10200 10320 10220 10360
rect 10260 10320 10280 10360
rect 10320 10320 10340 10360
rect 10380 10320 10400 10360
rect 8800 10080 9000 10100
rect 8800 10040 8820 10080
rect 8860 10040 8880 10080
rect 8920 10040 8940 10080
rect 8980 10040 9000 10080
rect 8800 10020 9000 10040
rect 8800 9980 8820 10020
rect 8860 9980 8880 10020
rect 8920 9980 8940 10020
rect 8980 9980 9000 10020
rect 8800 9960 9000 9980
rect 8800 9920 8820 9960
rect 8860 9920 8880 9960
rect 8920 9920 8940 9960
rect 8980 9920 9000 9960
rect 8800 580 9000 9920
rect 8800 540 8820 580
rect 8860 540 8880 580
rect 8920 540 8940 580
rect 8980 540 9000 580
rect 8800 520 9000 540
rect 8800 480 8820 520
rect 8860 480 8880 520
rect 8920 480 8940 520
rect 8980 480 9000 520
rect 8800 460 9000 480
rect 8800 420 8820 460
rect 8860 420 8880 460
rect 8920 420 8940 460
rect 8980 420 9000 460
rect 8800 400 9000 420
rect 7400 140 7420 180
rect 7460 140 7480 180
rect 7520 140 7540 180
rect 7580 140 7600 180
rect 7400 120 7600 140
rect 7400 80 7420 120
rect 7460 80 7480 120
rect 7520 80 7540 120
rect 7580 80 7600 120
rect 7400 60 7600 80
rect 7400 20 7420 60
rect 7460 20 7480 60
rect 7520 20 7540 60
rect 7580 20 7600 60
rect 7400 0 7600 20
rect 10200 180 10400 10320
rect 12000 10480 12200 10500
rect 12000 10440 12020 10480
rect 12060 10440 12080 10480
rect 12120 10440 12140 10480
rect 12180 10440 12200 10480
rect 12000 10420 12200 10440
rect 12000 10380 12020 10420
rect 12060 10380 12080 10420
rect 12120 10380 12140 10420
rect 12180 10380 12200 10420
rect 12000 10360 12200 10380
rect 12000 10320 12020 10360
rect 12060 10320 12080 10360
rect 12120 10320 12140 10360
rect 12180 10320 12200 10360
rect 11600 10080 11800 10100
rect 11600 10040 11620 10080
rect 11660 10040 11680 10080
rect 11720 10040 11740 10080
rect 11780 10040 11800 10080
rect 11600 10020 11800 10040
rect 11600 9980 11620 10020
rect 11660 9980 11680 10020
rect 11720 9980 11740 10020
rect 11780 9980 11800 10020
rect 11600 9960 11800 9980
rect 11600 9920 11620 9960
rect 11660 9920 11680 9960
rect 11720 9920 11740 9960
rect 11780 9920 11800 9960
rect 11600 580 11800 9920
rect 11600 540 11620 580
rect 11660 540 11680 580
rect 11720 540 11740 580
rect 11780 540 11800 580
rect 11600 520 11800 540
rect 11600 480 11620 520
rect 11660 480 11680 520
rect 11720 480 11740 520
rect 11780 480 11800 520
rect 11600 460 11800 480
rect 11600 420 11620 460
rect 11660 420 11680 460
rect 11720 420 11740 460
rect 11780 420 11800 460
rect 11600 400 11800 420
rect 10200 140 10220 180
rect 10260 140 10280 180
rect 10320 140 10340 180
rect 10380 140 10400 180
rect 10200 120 10400 140
rect 10200 80 10220 120
rect 10260 80 10280 120
rect 10320 80 10340 120
rect 10380 80 10400 120
rect 10200 60 10400 80
rect 10200 20 10220 60
rect 10260 20 10280 60
rect 10320 20 10340 60
rect 10380 20 10400 60
rect 10200 0 10400 20
rect 12000 180 12200 10320
rect 12000 140 12020 180
rect 12060 140 12080 180
rect 12120 140 12140 180
rect 12180 140 12200 180
rect 12000 120 12200 140
rect 12000 80 12020 120
rect 12060 80 12080 120
rect 12120 80 12140 120
rect 12180 80 12200 120
rect 12000 60 12200 80
rect 12000 20 12020 60
rect 12060 20 12080 60
rect 12120 20 12140 60
rect 12180 20 12200 60
rect 12000 0 12200 20
<< end >>
