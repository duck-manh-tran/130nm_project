magic
tech sky130A
magscale 1 2
timestamp 1624957691
<< psubdiff >>
rect 21600 6200 21602 6300
rect 21702 6200 21802 6300
rect 21902 6200 22000 6300
<< locali >>
rect 1229 12475 1398 12535
rect 476 12410 684 12420
rect 1688 12416 1732 12460
rect 476 12370 486 12410
rect 526 12370 684 12410
rect 476 12360 684 12370
rect 21600 6200 21602 6300
rect 21702 6280 21802 6300
rect 21902 6280 22000 6300
rect 21702 6220 21720 6280
rect 21780 6220 21802 6280
rect 21902 6220 21920 6280
rect 21980 6220 22000 6280
rect 21702 6200 21802 6220
rect 21902 6200 22000 6220
<< viali >>
rect 7220 14620 7280 14680
rect 7320 14620 7380 14680
rect 7420 14620 7480 14680
rect 7520 14620 7580 14680
rect 14420 14620 14480 14680
rect 14520 14620 14580 14680
rect 14620 14620 14680 14680
rect 14720 14620 14780 14680
rect 21620 14620 21680 14680
rect 21720 14620 21780 14680
rect 21820 14620 21880 14680
rect 21920 14620 21980 14680
rect 28820 14620 28880 14680
rect 28920 14620 28980 14680
rect 29020 14620 29080 14680
rect 29120 14620 29180 14680
rect 486 12370 526 12410
rect 7220 6220 7280 6280
rect 7320 6220 7380 6280
rect 7420 6220 7480 6280
rect 7520 6220 7580 6280
rect 14420 6220 14480 6280
rect 14520 6220 14580 6280
rect 14620 6220 14680 6280
rect 14720 6220 14780 6280
rect 21620 6220 21680 6280
rect 21720 6220 21780 6280
rect 21820 6220 21880 6280
rect 21920 6220 21980 6280
rect 28820 6220 28880 6280
rect 28920 6220 28980 6280
rect 29020 6220 29080 6280
rect 29120 6220 29180 6280
<< metal1 >>
rect 7200 14680 7600 14700
rect 7200 14620 7220 14680
rect 7286 14620 7298 14680
rect 7502 14620 7514 14680
rect 7580 14620 7600 14680
rect 7200 14600 7600 14620
rect 14400 14680 14800 14700
rect 14400 14620 14420 14680
rect 14486 14620 14498 14680
rect 14702 14620 14714 14680
rect 14780 14620 14800 14680
rect 14400 14600 14800 14620
rect 21600 14680 22000 14700
rect 21600 14620 21620 14680
rect 21686 14620 21698 14680
rect 21902 14620 21914 14680
rect 21980 14620 22000 14680
rect 21600 14600 22000 14620
rect 28800 14680 29200 14700
rect 28800 14620 28820 14680
rect 28886 14620 28898 14680
rect 29102 14620 29114 14680
rect 29180 14620 29200 14680
rect 28800 14600 29200 14620
rect 3102 13762 3974 13780
rect 3102 13702 3626 13762
rect 3686 13702 3698 13762
rect 3758 13702 3770 13762
rect 3830 13702 3842 13762
rect 3902 13702 3914 13762
rect 3102 13684 3974 13702
rect 10826 13762 11174 13780
rect 10886 13702 10898 13762
rect 10958 13702 10970 13762
rect 11030 13702 11042 13762
rect 11102 13702 11114 13762
rect 10826 13684 11174 13702
rect 18026 13762 18374 13780
rect 18086 13702 18098 13762
rect 18158 13702 18170 13762
rect 18230 13702 18242 13762
rect 18302 13702 18314 13762
rect 18026 13684 18374 13702
rect 25226 13762 25574 13780
rect 25286 13702 25298 13762
rect 25358 13702 25370 13762
rect 25430 13702 25442 13762
rect 25502 13702 25514 13762
rect 25226 13684 25574 13702
rect 32426 13762 32774 13780
rect 32486 13702 32498 13762
rect 32558 13702 32570 13762
rect 32630 13702 32642 13762
rect 32702 13702 32714 13762
rect 32426 13684 32774 13702
rect 9238 12852 9536 12980
rect 15150 12854 15448 12982
rect 21054 12852 21352 12980
rect 26946 12852 27244 12980
rect 2852 12674 4000 12692
rect 2852 12614 3626 12674
rect 3686 12614 3698 12674
rect 3758 12614 3770 12674
rect 3830 12614 3842 12674
rect 3902 12614 3914 12674
rect 3974 12614 4000 12674
rect 2852 12596 4000 12614
rect 474 12416 542 12420
rect 474 12364 480 12416
rect 532 12364 542 12416
rect 474 12360 542 12364
rect 0 12130 400 12148
rect 0 12070 26 12130
rect 86 12070 98 12130
rect 158 12070 170 12130
rect 230 12070 242 12130
rect 302 12070 314 12130
rect 374 12070 400 12130
rect 0 12052 400 12070
rect 35346 12130 36400 12148
rect 35346 12070 36026 12130
rect 36086 12070 36098 12130
rect 36158 12070 36170 12130
rect 36230 12070 36242 12130
rect 36302 12070 36314 12130
rect 36374 12070 36400 12130
rect 35346 12052 36400 12070
rect 2904 11586 3974 11604
rect 2904 11526 3626 11586
rect 3686 11526 3698 11586
rect 3758 11526 3770 11586
rect 3830 11526 3842 11586
rect 3902 11526 3914 11586
rect 2904 11508 3974 11526
rect 10826 11586 11174 11604
rect 10886 11526 10898 11586
rect 10958 11526 10970 11586
rect 11030 11526 11042 11586
rect 11102 11526 11114 11586
rect 10826 11508 11174 11526
rect 18026 11586 18374 11604
rect 18086 11526 18098 11586
rect 18158 11526 18170 11586
rect 18230 11526 18242 11586
rect 18302 11526 18314 11586
rect 18026 11508 18374 11526
rect 25226 11586 25574 11604
rect 25286 11526 25298 11586
rect 25358 11526 25370 11586
rect 25430 11526 25442 11586
rect 25502 11526 25514 11586
rect 25226 11508 25574 11526
rect 32426 11585 34192 11604
rect 32486 11525 32498 11585
rect 32558 11525 32570 11585
rect 32630 11525 32642 11585
rect 32702 11525 32714 11585
rect 32774 11525 34192 11585
rect 32426 11508 34192 11525
rect 32400 11507 32800 11508
rect 30904 10962 31422 11060
rect 0 9410 3974 9428
rect 0 9350 3626 9410
rect 3686 9350 3698 9410
rect 3758 9350 3770 9410
rect 3830 9350 3842 9410
rect 3902 9350 3914 9410
rect 0 9332 3974 9350
rect 10826 9410 11174 9428
rect 10886 9350 10898 9410
rect 10958 9350 10970 9410
rect 11030 9350 11042 9410
rect 11102 9350 11114 9410
rect 10826 9332 11174 9350
rect 18026 9410 18374 9428
rect 18086 9350 18098 9410
rect 18158 9350 18170 9410
rect 18230 9350 18242 9410
rect 18302 9350 18314 9410
rect 18026 9332 18374 9350
rect 25226 9410 25574 9428
rect 25286 9350 25298 9410
rect 25358 9350 25370 9410
rect 25430 9350 25442 9410
rect 25502 9350 25514 9410
rect 25226 9332 25574 9350
rect 32426 9410 35791 9428
rect 32486 9350 32498 9410
rect 32558 9350 32570 9410
rect 32630 9350 32642 9410
rect 32702 9350 32714 9410
rect 32774 9350 35791 9410
rect 32426 9332 35791 9350
rect 6046 7956 6344 8084
rect 11946 7954 12244 8082
rect 17858 7954 18156 8082
rect 23754 7954 24052 8082
rect 29670 7954 29968 8082
rect 0 7234 3974 7252
rect 0 7174 3626 7234
rect 3686 7174 3698 7234
rect 3758 7174 3770 7234
rect 3830 7174 3842 7234
rect 3902 7174 3914 7234
rect 0 7156 3974 7174
rect 10826 7234 11174 7252
rect 10886 7174 10898 7234
rect 10958 7174 10970 7234
rect 11030 7174 11042 7234
rect 11102 7174 11114 7234
rect 10826 7156 11174 7174
rect 25226 7234 25574 7252
rect 25286 7174 25298 7234
rect 25358 7174 25370 7234
rect 25430 7174 25442 7234
rect 25502 7174 25514 7234
rect 25226 7156 25574 7174
rect 32426 7234 35790 7252
rect 32486 7174 32498 7234
rect 32558 7174 32570 7234
rect 32630 7174 32642 7234
rect 32702 7174 32714 7234
rect 32774 7174 35790 7234
rect 32426 7156 35790 7174
rect 7200 6280 7600 6300
rect 7200 6220 7220 6280
rect 7286 6220 7298 6280
rect 7502 6220 7514 6280
rect 7580 6220 7600 6280
rect 7200 6212 7600 6220
rect 14400 6280 14800 6300
rect 14400 6220 14420 6280
rect 14486 6220 14498 6280
rect 14702 6220 14714 6280
rect 14780 6220 14800 6280
rect 7200 6200 7528 6212
rect 14400 6200 14800 6220
rect 21600 6280 22000 6300
rect 21600 6220 21620 6280
rect 21686 6220 21698 6280
rect 21902 6220 21914 6280
rect 21980 6220 22000 6280
rect 21600 6200 22000 6220
rect 28800 6280 29200 6300
rect 28800 6220 28820 6280
rect 28886 6220 28898 6280
rect 29102 6220 29114 6280
rect 29180 6220 29200 6280
rect 28800 6200 29200 6220
<< via1 >>
rect 7226 14620 7280 14680
rect 7280 14620 7286 14680
rect 7298 14620 7320 14680
rect 7320 14620 7358 14680
rect 7370 14620 7380 14680
rect 7380 14620 7420 14680
rect 7420 14620 7430 14680
rect 7442 14620 7480 14680
rect 7480 14620 7502 14680
rect 7514 14620 7520 14680
rect 7520 14620 7574 14680
rect 14426 14620 14480 14680
rect 14480 14620 14486 14680
rect 14498 14620 14520 14680
rect 14520 14620 14558 14680
rect 14570 14620 14580 14680
rect 14580 14620 14620 14680
rect 14620 14620 14630 14680
rect 14642 14620 14680 14680
rect 14680 14620 14702 14680
rect 14714 14620 14720 14680
rect 14720 14620 14774 14680
rect 21626 14620 21680 14680
rect 21680 14620 21686 14680
rect 21698 14620 21720 14680
rect 21720 14620 21758 14680
rect 21770 14620 21780 14680
rect 21780 14620 21820 14680
rect 21820 14620 21830 14680
rect 21842 14620 21880 14680
rect 21880 14620 21902 14680
rect 21914 14620 21920 14680
rect 21920 14620 21974 14680
rect 28826 14620 28880 14680
rect 28880 14620 28886 14680
rect 28898 14620 28920 14680
rect 28920 14620 28958 14680
rect 28970 14620 28980 14680
rect 28980 14620 29020 14680
rect 29020 14620 29030 14680
rect 29042 14620 29080 14680
rect 29080 14620 29102 14680
rect 29114 14620 29120 14680
rect 29120 14620 29174 14680
rect 3626 13702 3686 13762
rect 3698 13702 3758 13762
rect 3770 13702 3830 13762
rect 3842 13702 3902 13762
rect 3914 13702 3974 13762
rect 10826 13702 10886 13762
rect 10898 13702 10958 13762
rect 10970 13702 11030 13762
rect 11042 13702 11102 13762
rect 11114 13702 11174 13762
rect 18026 13702 18086 13762
rect 18098 13702 18158 13762
rect 18170 13702 18230 13762
rect 18242 13702 18302 13762
rect 18314 13702 18374 13762
rect 25226 13702 25286 13762
rect 25298 13702 25358 13762
rect 25370 13702 25430 13762
rect 25442 13702 25502 13762
rect 25514 13702 25574 13762
rect 32426 13702 32486 13762
rect 32498 13702 32558 13762
rect 32570 13702 32630 13762
rect 32642 13702 32702 13762
rect 32714 13702 32774 13762
rect 3626 12614 3686 12674
rect 3698 12614 3758 12674
rect 3770 12614 3830 12674
rect 3842 12614 3902 12674
rect 3914 12614 3974 12674
rect 480 12410 532 12416
rect 480 12370 486 12410
rect 486 12370 526 12410
rect 526 12370 532 12410
rect 480 12364 532 12370
rect 9258 12340 9322 12404
rect 9354 12342 9418 12406
rect 15146 12340 15210 12404
rect 15242 12342 15306 12406
rect 21034 12340 21098 12404
rect 21130 12342 21194 12406
rect 26922 12340 26986 12404
rect 27018 12342 27082 12406
rect 26 12070 86 12130
rect 98 12070 158 12130
rect 170 12070 230 12130
rect 242 12070 302 12130
rect 314 12070 374 12130
rect 36026 12070 36086 12130
rect 36098 12070 36158 12130
rect 36170 12070 36230 12130
rect 36242 12070 36302 12130
rect 36314 12070 36374 12130
rect 3626 11526 3686 11586
rect 3698 11526 3758 11586
rect 3770 11526 3830 11586
rect 3842 11526 3902 11586
rect 3914 11526 3974 11586
rect 10826 11526 10886 11586
rect 10898 11526 10958 11586
rect 10970 11526 11030 11586
rect 11042 11526 11102 11586
rect 11114 11526 11174 11586
rect 18026 11526 18086 11586
rect 18098 11526 18158 11586
rect 18170 11526 18230 11586
rect 18242 11526 18302 11586
rect 18314 11526 18374 11586
rect 25226 11526 25286 11586
rect 25298 11526 25358 11586
rect 25370 11526 25430 11586
rect 25442 11526 25502 11586
rect 25514 11526 25574 11586
rect 32426 11525 32486 11585
rect 32498 11525 32558 11585
rect 32570 11525 32630 11585
rect 32642 11525 32702 11585
rect 32714 11525 32774 11585
rect 3626 9350 3686 9410
rect 3698 9350 3758 9410
rect 3770 9350 3830 9410
rect 3842 9350 3902 9410
rect 3914 9350 3974 9410
rect 10826 9350 10886 9410
rect 10898 9350 10958 9410
rect 10970 9350 11030 9410
rect 11042 9350 11102 9410
rect 11114 9350 11174 9410
rect 18026 9350 18086 9410
rect 18098 9350 18158 9410
rect 18170 9350 18230 9410
rect 18242 9350 18302 9410
rect 18314 9350 18374 9410
rect 25226 9350 25286 9410
rect 25298 9350 25358 9410
rect 25370 9350 25430 9410
rect 25442 9350 25502 9410
rect 25514 9350 25574 9410
rect 32426 9350 32486 9410
rect 32498 9350 32558 9410
rect 32570 9350 32630 9410
rect 32642 9350 32702 9410
rect 32714 9350 32774 9410
rect 6130 8524 6194 8588
rect 6226 8526 6290 8590
rect 12018 8524 12082 8588
rect 12114 8526 12178 8590
rect 17906 8524 17970 8588
rect 18002 8526 18066 8590
rect 23886 8524 23950 8588
rect 23982 8526 24046 8590
rect 29774 8524 29838 8588
rect 29870 8526 29934 8590
rect 3626 7174 3686 7234
rect 3698 7174 3758 7234
rect 3770 7174 3830 7234
rect 3842 7174 3902 7234
rect 3914 7174 3974 7234
rect 10826 7174 10886 7234
rect 10898 7174 10958 7234
rect 10970 7174 11030 7234
rect 11042 7174 11102 7234
rect 11114 7174 11174 7234
rect 25226 7174 25286 7234
rect 25298 7174 25358 7234
rect 25370 7174 25430 7234
rect 25442 7174 25502 7234
rect 25514 7174 25574 7234
rect 32426 7174 32486 7234
rect 32498 7174 32558 7234
rect 32570 7174 32630 7234
rect 32642 7174 32702 7234
rect 32714 7174 32774 7234
rect 7226 6220 7280 6280
rect 7280 6220 7286 6280
rect 7298 6220 7320 6280
rect 7320 6220 7358 6280
rect 7370 6220 7380 6280
rect 7380 6220 7420 6280
rect 7420 6220 7430 6280
rect 7442 6220 7480 6280
rect 7480 6220 7502 6280
rect 7514 6220 7520 6280
rect 7520 6220 7574 6280
rect 14426 6220 14480 6280
rect 14480 6220 14486 6280
rect 14498 6220 14520 6280
rect 14520 6220 14558 6280
rect 14570 6220 14580 6280
rect 14580 6220 14620 6280
rect 14620 6220 14630 6280
rect 14642 6220 14680 6280
rect 14680 6220 14702 6280
rect 14714 6220 14720 6280
rect 14720 6220 14774 6280
rect 21626 6220 21680 6280
rect 21680 6220 21686 6280
rect 21698 6220 21720 6280
rect 21720 6220 21758 6280
rect 21770 6220 21780 6280
rect 21780 6220 21820 6280
rect 21820 6220 21830 6280
rect 21842 6220 21880 6280
rect 21880 6220 21902 6280
rect 21914 6220 21920 6280
rect 21920 6220 21974 6280
rect 28826 6220 28880 6280
rect 28880 6220 28886 6280
rect 28898 6220 28920 6280
rect 28920 6220 28958 6280
rect 28970 6220 28980 6280
rect 28980 6220 29020 6280
rect 29020 6220 29030 6280
rect 29042 6220 29080 6280
rect 29080 6220 29102 6280
rect 29114 6220 29120 6280
rect 29120 6220 29174 6280
<< metal2 >>
rect 7200 14682 7600 14700
rect 7200 14680 7236 14682
rect 7300 14680 7324 14682
rect 7388 14680 7412 14682
rect 7476 14680 7500 14682
rect 7564 14680 7600 14682
rect 7200 14620 7226 14680
rect 7574 14620 7600 14680
rect 7200 14618 7236 14620
rect 7300 14618 7324 14620
rect 7388 14618 7412 14620
rect 7476 14618 7500 14620
rect 7564 14618 7600 14620
rect 7200 14600 7600 14618
rect 14400 14682 14800 14700
rect 14400 14680 14436 14682
rect 14500 14680 14524 14682
rect 14588 14680 14612 14682
rect 14676 14680 14700 14682
rect 14764 14680 14800 14682
rect 14400 14620 14426 14680
rect 14774 14620 14800 14680
rect 14400 14618 14436 14620
rect 14500 14618 14524 14620
rect 14588 14618 14612 14620
rect 14676 14618 14700 14620
rect 14764 14618 14800 14620
rect 14400 14600 14800 14618
rect 21600 14682 22000 14700
rect 21600 14680 21636 14682
rect 21700 14680 21724 14682
rect 21788 14680 21812 14682
rect 21876 14680 21900 14682
rect 21964 14680 22000 14682
rect 21600 14620 21626 14680
rect 21974 14620 22000 14680
rect 21600 14618 21636 14620
rect 21700 14618 21724 14620
rect 21788 14618 21812 14620
rect 21876 14618 21900 14620
rect 21964 14618 22000 14620
rect 21600 14600 22000 14618
rect 28800 14682 29200 14700
rect 28800 14680 28836 14682
rect 28900 14680 28924 14682
rect 28988 14680 29012 14682
rect 29076 14680 29100 14682
rect 29164 14680 29200 14682
rect 28800 14620 28826 14680
rect 29174 14620 29200 14680
rect 28800 14618 28836 14620
rect 28900 14618 28924 14620
rect 28988 14618 29012 14620
rect 29076 14618 29100 14620
rect 29164 14618 29200 14620
rect 28800 14600 29200 14618
rect 3600 13764 4000 13780
rect 3600 13762 3636 13764
rect 3700 13762 3724 13764
rect 3788 13762 3812 13764
rect 3876 13762 3900 13764
rect 3964 13762 4000 13764
rect 3600 13702 3626 13762
rect 3974 13702 4000 13762
rect 3600 13700 3636 13702
rect 3700 13700 3724 13702
rect 3788 13700 3812 13702
rect 3876 13700 3900 13702
rect 3964 13700 4000 13702
rect 3600 13684 4000 13700
rect 10800 13764 11200 13780
rect 10800 13762 10836 13764
rect 10900 13762 10924 13764
rect 10988 13762 11012 13764
rect 11076 13762 11100 13764
rect 11164 13762 11200 13764
rect 10800 13702 10826 13762
rect 11174 13702 11200 13762
rect 10800 13700 10836 13702
rect 10900 13700 10924 13702
rect 10988 13700 11012 13702
rect 11076 13700 11100 13702
rect 11164 13700 11200 13702
rect 10800 13684 11200 13700
rect 18000 13764 18400 13780
rect 18000 13762 18036 13764
rect 18100 13762 18124 13764
rect 18188 13762 18212 13764
rect 18276 13762 18300 13764
rect 18364 13762 18400 13764
rect 18000 13702 18026 13762
rect 18374 13702 18400 13762
rect 18000 13700 18036 13702
rect 18100 13700 18124 13702
rect 18188 13700 18212 13702
rect 18276 13700 18300 13702
rect 18364 13700 18400 13702
rect 18000 13684 18400 13700
rect 25200 13764 25600 13780
rect 25200 13762 25236 13764
rect 25300 13762 25324 13764
rect 25388 13762 25412 13764
rect 25476 13762 25500 13764
rect 25564 13762 25600 13764
rect 25200 13702 25226 13762
rect 25574 13702 25600 13762
rect 25200 13700 25236 13702
rect 25300 13700 25324 13702
rect 25388 13700 25412 13702
rect 25476 13700 25500 13702
rect 25564 13700 25600 13702
rect 25200 13684 25600 13700
rect 32400 13764 32800 13780
rect 32400 13762 32436 13764
rect 32500 13762 32524 13764
rect 32588 13762 32612 13764
rect 32676 13762 32700 13764
rect 32764 13762 32800 13764
rect 32400 13702 32426 13762
rect 32774 13702 32800 13762
rect 32400 13700 32436 13702
rect 32500 13700 32524 13702
rect 32588 13700 32612 13702
rect 32676 13700 32700 13702
rect 32764 13700 32800 13702
rect 32400 13684 32800 13700
rect 3600 12676 4000 12692
rect 3600 12674 3636 12676
rect 3700 12674 3724 12676
rect 3788 12674 3812 12676
rect 3876 12674 3900 12676
rect 3964 12674 4000 12676
rect 3600 12614 3626 12674
rect 3974 12614 4000 12674
rect 3600 12612 3636 12614
rect 3700 12612 3724 12614
rect 3788 12612 3812 12614
rect 3876 12612 3900 12614
rect 3964 12612 4000 12614
rect 3600 12596 4000 12612
rect 466 12360 476 12420
rect 536 12360 546 12420
rect 9246 12406 9430 12418
rect 9246 12404 9354 12406
rect 9246 12340 9258 12404
rect 9322 12342 9354 12404
rect 9418 12342 9430 12406
rect 9322 12340 9430 12342
rect 9246 12326 9430 12340
rect 15134 12406 15318 12418
rect 15134 12404 15242 12406
rect 15134 12340 15146 12404
rect 15210 12342 15242 12404
rect 15306 12342 15318 12406
rect 15210 12340 15318 12342
rect 15134 12326 15318 12340
rect 21022 12406 21206 12418
rect 21022 12404 21130 12406
rect 21022 12340 21034 12404
rect 21098 12342 21130 12404
rect 21194 12342 21206 12406
rect 21098 12340 21206 12342
rect 21022 12326 21206 12340
rect 26910 12406 27094 12418
rect 26910 12404 27018 12406
rect 26910 12340 26922 12404
rect 26986 12342 27018 12404
rect 27082 12342 27094 12406
rect 26986 12340 27094 12342
rect 26910 12326 27094 12340
rect 0 12132 400 12148
rect 0 12130 36 12132
rect 100 12130 124 12132
rect 188 12130 212 12132
rect 276 12130 300 12132
rect 364 12130 400 12132
rect 0 12070 26 12130
rect 374 12070 400 12130
rect 0 12068 36 12070
rect 100 12068 124 12070
rect 188 12068 212 12070
rect 276 12068 300 12070
rect 364 12068 400 12070
rect 0 12052 400 12068
rect 36000 12132 36400 12148
rect 36000 12130 36036 12132
rect 36100 12130 36124 12132
rect 36188 12130 36212 12132
rect 36276 12130 36300 12132
rect 36364 12130 36400 12132
rect 36000 12070 36026 12130
rect 36374 12070 36400 12130
rect 36000 12068 36036 12070
rect 36100 12068 36124 12070
rect 36188 12068 36212 12070
rect 36276 12068 36300 12070
rect 36364 12068 36400 12070
rect 36000 12052 36400 12068
rect 35852 11738 36702 11898
rect 3600 11588 4000 11604
rect 3600 11586 3636 11588
rect 3700 11586 3724 11588
rect 3788 11586 3812 11588
rect 3876 11586 3900 11588
rect 3964 11586 4000 11588
rect 3600 11526 3626 11586
rect 3974 11526 4000 11586
rect 3600 11524 3636 11526
rect 3700 11524 3724 11526
rect 3788 11524 3812 11526
rect 3876 11524 3900 11526
rect 3964 11524 4000 11526
rect 3600 11508 4000 11524
rect 10800 11588 11200 11604
rect 10800 11586 10836 11588
rect 10900 11586 10924 11588
rect 10988 11586 11012 11588
rect 11076 11586 11100 11588
rect 11164 11586 11200 11588
rect 10800 11526 10826 11586
rect 11174 11526 11200 11586
rect 10800 11524 10836 11526
rect 10900 11524 10924 11526
rect 10988 11524 11012 11526
rect 11076 11524 11100 11526
rect 11164 11524 11200 11526
rect 10800 11508 11200 11524
rect 18000 11588 18400 11604
rect 18000 11586 18036 11588
rect 18100 11586 18124 11588
rect 18188 11586 18212 11588
rect 18276 11586 18300 11588
rect 18364 11586 18400 11588
rect 18000 11526 18026 11586
rect 18374 11526 18400 11586
rect 18000 11524 18036 11526
rect 18100 11524 18124 11526
rect 18188 11524 18212 11526
rect 18276 11524 18300 11526
rect 18364 11524 18400 11526
rect 18000 11508 18400 11524
rect 25200 11588 25600 11604
rect 25200 11586 25236 11588
rect 25300 11586 25324 11588
rect 25388 11586 25412 11588
rect 25476 11586 25500 11588
rect 25564 11586 25600 11588
rect 25200 11526 25226 11586
rect 25574 11526 25600 11586
rect 25200 11524 25236 11526
rect 25300 11524 25324 11526
rect 25388 11524 25412 11526
rect 25476 11524 25500 11526
rect 25564 11524 25600 11526
rect 25200 11508 25600 11524
rect 32400 11587 32800 11604
rect 32400 11585 32436 11587
rect 32500 11585 32524 11587
rect 32588 11585 32612 11587
rect 32676 11585 32700 11587
rect 32764 11585 32800 11587
rect 32400 11525 32426 11585
rect 32774 11525 32800 11585
rect 32400 11523 32436 11525
rect 32500 11523 32524 11525
rect 32588 11523 32612 11525
rect 32676 11523 32700 11525
rect 32764 11523 32800 11525
rect 32400 11507 32800 11523
rect 702 10532 1018 10670
rect 34266 10048 34582 10186
rect 3600 9412 4000 9428
rect 3600 9410 3636 9412
rect 3700 9410 3724 9412
rect 3788 9410 3812 9412
rect 3876 9410 3900 9412
rect 3964 9410 4000 9412
rect 3600 9350 3626 9410
rect 3974 9350 4000 9410
rect 3600 9348 3636 9350
rect 3700 9348 3724 9350
rect 3788 9348 3812 9350
rect 3876 9348 3900 9350
rect 3964 9348 4000 9350
rect 3600 9332 4000 9348
rect 10800 9412 11200 9428
rect 10800 9410 10836 9412
rect 10900 9410 10924 9412
rect 10988 9410 11012 9412
rect 11076 9410 11100 9412
rect 11164 9410 11200 9412
rect 10800 9350 10826 9410
rect 11174 9350 11200 9410
rect 10800 9348 10836 9350
rect 10900 9348 10924 9350
rect 10988 9348 11012 9350
rect 11076 9348 11100 9350
rect 11164 9348 11200 9350
rect 10800 9332 11200 9348
rect 18000 9412 18400 9428
rect 18000 9410 18036 9412
rect 18100 9410 18124 9412
rect 18188 9410 18212 9412
rect 18276 9410 18300 9412
rect 18364 9410 18400 9412
rect 18000 9350 18026 9410
rect 18374 9350 18400 9410
rect 18000 9348 18036 9350
rect 18100 9348 18124 9350
rect 18188 9348 18212 9350
rect 18276 9348 18300 9350
rect 18364 9348 18400 9350
rect 18000 9332 18400 9348
rect 25200 9412 25600 9428
rect 25200 9410 25236 9412
rect 25300 9410 25324 9412
rect 25388 9410 25412 9412
rect 25476 9410 25500 9412
rect 25564 9410 25600 9412
rect 25200 9350 25226 9410
rect 25574 9350 25600 9410
rect 25200 9348 25236 9350
rect 25300 9348 25324 9350
rect 25388 9348 25412 9350
rect 25476 9348 25500 9350
rect 25564 9348 25600 9350
rect 25200 9332 25600 9348
rect 32400 9412 32800 9428
rect 32400 9410 32436 9412
rect 32500 9410 32524 9412
rect 32588 9410 32612 9412
rect 32676 9410 32700 9412
rect 32764 9410 32800 9412
rect 32400 9350 32426 9410
rect 32774 9350 32800 9410
rect 32400 9348 32436 9350
rect 32500 9348 32524 9350
rect 32588 9348 32612 9350
rect 32676 9348 32700 9350
rect 32764 9348 32800 9350
rect 32400 9332 32800 9348
rect 1228 8510 1412 8602
rect 6118 8590 6302 8602
rect 6118 8588 6226 8590
rect 6118 8524 6130 8588
rect 6194 8526 6226 8588
rect 6290 8526 6302 8590
rect 6194 8524 6302 8526
rect 6118 8510 6302 8524
rect 12006 8590 12190 8602
rect 12006 8588 12114 8590
rect 12006 8524 12018 8588
rect 12082 8526 12114 8588
rect 12178 8526 12190 8590
rect 12082 8524 12190 8526
rect 12006 8510 12190 8524
rect 17894 8590 18078 8602
rect 17894 8588 18002 8590
rect 17894 8524 17906 8588
rect 17970 8526 18002 8588
rect 18066 8526 18078 8590
rect 17970 8524 18078 8526
rect 17894 8510 18078 8524
rect 23874 8590 24058 8602
rect 23874 8588 23982 8590
rect 23874 8524 23886 8588
rect 23950 8526 23982 8588
rect 24046 8526 24058 8590
rect 23950 8524 24058 8526
rect 23874 8510 24058 8524
rect 29762 8590 29946 8602
rect 29762 8588 29870 8590
rect 29762 8524 29774 8588
rect 29838 8526 29870 8588
rect 29934 8526 29946 8590
rect 29838 8524 29946 8526
rect 29762 8510 29946 8524
rect 33166 8510 33350 8602
rect 3600 7236 4000 7252
rect 3600 7234 3636 7236
rect 3700 7234 3724 7236
rect 3788 7234 3812 7236
rect 3876 7234 3900 7236
rect 3964 7234 4000 7236
rect 3600 7174 3626 7234
rect 3974 7174 4000 7234
rect 3600 7172 3636 7174
rect 3700 7172 3724 7174
rect 3788 7172 3812 7174
rect 3876 7172 3900 7174
rect 3964 7172 4000 7174
rect 3600 7156 4000 7172
rect 10800 7236 11200 7252
rect 10800 7234 10836 7236
rect 10900 7234 10924 7236
rect 10988 7234 11012 7236
rect 11076 7234 11100 7236
rect 11164 7234 11200 7236
rect 10800 7174 10826 7234
rect 11174 7174 11200 7234
rect 10800 7172 10836 7174
rect 10900 7172 10924 7174
rect 10988 7172 11012 7174
rect 11076 7172 11100 7174
rect 11164 7172 11200 7174
rect 10800 7156 11200 7172
rect 25200 7236 25600 7252
rect 25200 7234 25236 7236
rect 25300 7234 25324 7236
rect 25388 7234 25412 7236
rect 25476 7234 25500 7236
rect 25564 7234 25600 7236
rect 25200 7174 25226 7234
rect 25574 7174 25600 7234
rect 25200 7172 25236 7174
rect 25300 7172 25324 7174
rect 25388 7172 25412 7174
rect 25476 7172 25500 7174
rect 25564 7172 25600 7174
rect 25200 7156 25600 7172
rect 32400 7236 32800 7252
rect 32400 7234 32436 7236
rect 32500 7234 32524 7236
rect 32588 7234 32612 7236
rect 32676 7234 32700 7236
rect 32764 7234 32800 7236
rect 32400 7174 32426 7234
rect 32774 7174 32800 7234
rect 32400 7172 32436 7174
rect 32500 7172 32524 7174
rect 32588 7172 32612 7174
rect 32676 7172 32700 7174
rect 32764 7172 32800 7174
rect 32400 7156 32800 7172
rect 7200 6282 7600 6300
rect 7200 6280 7236 6282
rect 7300 6280 7324 6282
rect 7388 6280 7412 6282
rect 7476 6280 7500 6282
rect 7564 6280 7600 6282
rect 7200 6220 7226 6280
rect 7574 6220 7600 6280
rect 7200 6218 7236 6220
rect 7300 6218 7324 6220
rect 7388 6218 7412 6220
rect 7476 6218 7500 6220
rect 7564 6218 7600 6220
rect 7200 6212 7600 6218
rect 14400 6282 14800 6300
rect 14400 6280 14436 6282
rect 14500 6280 14524 6282
rect 14588 6280 14612 6282
rect 14676 6280 14700 6282
rect 14764 6280 14800 6282
rect 14400 6220 14426 6280
rect 14774 6220 14800 6280
rect 14400 6218 14436 6220
rect 14500 6218 14524 6220
rect 14588 6218 14612 6220
rect 14676 6218 14700 6220
rect 14764 6218 14800 6220
rect 7200 6200 7528 6212
rect 14400 6200 14800 6218
rect 21600 6282 22000 6300
rect 21600 6280 21636 6282
rect 21700 6280 21724 6282
rect 21788 6280 21812 6282
rect 21876 6280 21900 6282
rect 21964 6280 22000 6282
rect 21600 6220 21626 6280
rect 21974 6220 22000 6280
rect 21600 6218 21636 6220
rect 21700 6218 21724 6220
rect 21788 6218 21812 6220
rect 21876 6218 21900 6220
rect 21964 6218 22000 6220
rect 21600 6200 22000 6218
rect 28800 6282 29200 6300
rect 28800 6280 28836 6282
rect 28900 6280 28924 6282
rect 28988 6280 29012 6282
rect 29076 6280 29100 6282
rect 29164 6280 29200 6282
rect 28800 6220 28826 6280
rect 29174 6220 29200 6280
rect 28800 6218 28836 6220
rect 28900 6218 28924 6220
rect 28988 6218 29012 6220
rect 29076 6218 29100 6220
rect 29164 6218 29200 6220
rect 28800 6200 29200 6218
<< via2 >>
rect 7236 14680 7300 14682
rect 7324 14680 7388 14682
rect 7412 14680 7476 14682
rect 7500 14680 7564 14682
rect 7236 14620 7286 14680
rect 7286 14620 7298 14680
rect 7298 14620 7300 14680
rect 7324 14620 7358 14680
rect 7358 14620 7370 14680
rect 7370 14620 7388 14680
rect 7412 14620 7430 14680
rect 7430 14620 7442 14680
rect 7442 14620 7476 14680
rect 7500 14620 7502 14680
rect 7502 14620 7514 14680
rect 7514 14620 7564 14680
rect 7236 14618 7300 14620
rect 7324 14618 7388 14620
rect 7412 14618 7476 14620
rect 7500 14618 7564 14620
rect 14436 14680 14500 14682
rect 14524 14680 14588 14682
rect 14612 14680 14676 14682
rect 14700 14680 14764 14682
rect 14436 14620 14486 14680
rect 14486 14620 14498 14680
rect 14498 14620 14500 14680
rect 14524 14620 14558 14680
rect 14558 14620 14570 14680
rect 14570 14620 14588 14680
rect 14612 14620 14630 14680
rect 14630 14620 14642 14680
rect 14642 14620 14676 14680
rect 14700 14620 14702 14680
rect 14702 14620 14714 14680
rect 14714 14620 14764 14680
rect 14436 14618 14500 14620
rect 14524 14618 14588 14620
rect 14612 14618 14676 14620
rect 14700 14618 14764 14620
rect 21636 14680 21700 14682
rect 21724 14680 21788 14682
rect 21812 14680 21876 14682
rect 21900 14680 21964 14682
rect 21636 14620 21686 14680
rect 21686 14620 21698 14680
rect 21698 14620 21700 14680
rect 21724 14620 21758 14680
rect 21758 14620 21770 14680
rect 21770 14620 21788 14680
rect 21812 14620 21830 14680
rect 21830 14620 21842 14680
rect 21842 14620 21876 14680
rect 21900 14620 21902 14680
rect 21902 14620 21914 14680
rect 21914 14620 21964 14680
rect 21636 14618 21700 14620
rect 21724 14618 21788 14620
rect 21812 14618 21876 14620
rect 21900 14618 21964 14620
rect 28836 14680 28900 14682
rect 28924 14680 28988 14682
rect 29012 14680 29076 14682
rect 29100 14680 29164 14682
rect 28836 14620 28886 14680
rect 28886 14620 28898 14680
rect 28898 14620 28900 14680
rect 28924 14620 28958 14680
rect 28958 14620 28970 14680
rect 28970 14620 28988 14680
rect 29012 14620 29030 14680
rect 29030 14620 29042 14680
rect 29042 14620 29076 14680
rect 29100 14620 29102 14680
rect 29102 14620 29114 14680
rect 29114 14620 29164 14680
rect 28836 14618 28900 14620
rect 28924 14618 28988 14620
rect 29012 14618 29076 14620
rect 29100 14618 29164 14620
rect 3636 13762 3700 13764
rect 3724 13762 3788 13764
rect 3812 13762 3876 13764
rect 3900 13762 3964 13764
rect 3636 13702 3686 13762
rect 3686 13702 3698 13762
rect 3698 13702 3700 13762
rect 3724 13702 3758 13762
rect 3758 13702 3770 13762
rect 3770 13702 3788 13762
rect 3812 13702 3830 13762
rect 3830 13702 3842 13762
rect 3842 13702 3876 13762
rect 3900 13702 3902 13762
rect 3902 13702 3914 13762
rect 3914 13702 3964 13762
rect 3636 13700 3700 13702
rect 3724 13700 3788 13702
rect 3812 13700 3876 13702
rect 3900 13700 3964 13702
rect 10836 13762 10900 13764
rect 10924 13762 10988 13764
rect 11012 13762 11076 13764
rect 11100 13762 11164 13764
rect 10836 13702 10886 13762
rect 10886 13702 10898 13762
rect 10898 13702 10900 13762
rect 10924 13702 10958 13762
rect 10958 13702 10970 13762
rect 10970 13702 10988 13762
rect 11012 13702 11030 13762
rect 11030 13702 11042 13762
rect 11042 13702 11076 13762
rect 11100 13702 11102 13762
rect 11102 13702 11114 13762
rect 11114 13702 11164 13762
rect 10836 13700 10900 13702
rect 10924 13700 10988 13702
rect 11012 13700 11076 13702
rect 11100 13700 11164 13702
rect 18036 13762 18100 13764
rect 18124 13762 18188 13764
rect 18212 13762 18276 13764
rect 18300 13762 18364 13764
rect 18036 13702 18086 13762
rect 18086 13702 18098 13762
rect 18098 13702 18100 13762
rect 18124 13702 18158 13762
rect 18158 13702 18170 13762
rect 18170 13702 18188 13762
rect 18212 13702 18230 13762
rect 18230 13702 18242 13762
rect 18242 13702 18276 13762
rect 18300 13702 18302 13762
rect 18302 13702 18314 13762
rect 18314 13702 18364 13762
rect 18036 13700 18100 13702
rect 18124 13700 18188 13702
rect 18212 13700 18276 13702
rect 18300 13700 18364 13702
rect 25236 13762 25300 13764
rect 25324 13762 25388 13764
rect 25412 13762 25476 13764
rect 25500 13762 25564 13764
rect 25236 13702 25286 13762
rect 25286 13702 25298 13762
rect 25298 13702 25300 13762
rect 25324 13702 25358 13762
rect 25358 13702 25370 13762
rect 25370 13702 25388 13762
rect 25412 13702 25430 13762
rect 25430 13702 25442 13762
rect 25442 13702 25476 13762
rect 25500 13702 25502 13762
rect 25502 13702 25514 13762
rect 25514 13702 25564 13762
rect 25236 13700 25300 13702
rect 25324 13700 25388 13702
rect 25412 13700 25476 13702
rect 25500 13700 25564 13702
rect 32436 13762 32500 13764
rect 32524 13762 32588 13764
rect 32612 13762 32676 13764
rect 32700 13762 32764 13764
rect 32436 13702 32486 13762
rect 32486 13702 32498 13762
rect 32498 13702 32500 13762
rect 32524 13702 32558 13762
rect 32558 13702 32570 13762
rect 32570 13702 32588 13762
rect 32612 13702 32630 13762
rect 32630 13702 32642 13762
rect 32642 13702 32676 13762
rect 32700 13702 32702 13762
rect 32702 13702 32714 13762
rect 32714 13702 32764 13762
rect 32436 13700 32500 13702
rect 32524 13700 32588 13702
rect 32612 13700 32676 13702
rect 32700 13700 32764 13702
rect 3636 12674 3700 12676
rect 3724 12674 3788 12676
rect 3812 12674 3876 12676
rect 3900 12674 3964 12676
rect 3636 12614 3686 12674
rect 3686 12614 3698 12674
rect 3698 12614 3700 12674
rect 3724 12614 3758 12674
rect 3758 12614 3770 12674
rect 3770 12614 3788 12674
rect 3812 12614 3830 12674
rect 3830 12614 3842 12674
rect 3842 12614 3876 12674
rect 3900 12614 3902 12674
rect 3902 12614 3914 12674
rect 3914 12614 3964 12674
rect 3636 12612 3700 12614
rect 3724 12612 3788 12614
rect 3812 12612 3876 12614
rect 3900 12612 3964 12614
rect 476 12416 536 12420
rect 476 12364 480 12416
rect 480 12364 532 12416
rect 532 12364 536 12416
rect 476 12360 536 12364
rect 36 12130 100 12132
rect 124 12130 188 12132
rect 212 12130 276 12132
rect 300 12130 364 12132
rect 36 12070 86 12130
rect 86 12070 98 12130
rect 98 12070 100 12130
rect 124 12070 158 12130
rect 158 12070 170 12130
rect 170 12070 188 12130
rect 212 12070 230 12130
rect 230 12070 242 12130
rect 242 12070 276 12130
rect 300 12070 302 12130
rect 302 12070 314 12130
rect 314 12070 364 12130
rect 36 12068 100 12070
rect 124 12068 188 12070
rect 212 12068 276 12070
rect 300 12068 364 12070
rect 36036 12130 36100 12132
rect 36124 12130 36188 12132
rect 36212 12130 36276 12132
rect 36300 12130 36364 12132
rect 36036 12070 36086 12130
rect 36086 12070 36098 12130
rect 36098 12070 36100 12130
rect 36124 12070 36158 12130
rect 36158 12070 36170 12130
rect 36170 12070 36188 12130
rect 36212 12070 36230 12130
rect 36230 12070 36242 12130
rect 36242 12070 36276 12130
rect 36300 12070 36302 12130
rect 36302 12070 36314 12130
rect 36314 12070 36364 12130
rect 36036 12068 36100 12070
rect 36124 12068 36188 12070
rect 36212 12068 36276 12070
rect 36300 12068 36364 12070
rect 3636 11586 3700 11588
rect 3724 11586 3788 11588
rect 3812 11586 3876 11588
rect 3900 11586 3964 11588
rect 3636 11526 3686 11586
rect 3686 11526 3698 11586
rect 3698 11526 3700 11586
rect 3724 11526 3758 11586
rect 3758 11526 3770 11586
rect 3770 11526 3788 11586
rect 3812 11526 3830 11586
rect 3830 11526 3842 11586
rect 3842 11526 3876 11586
rect 3900 11526 3902 11586
rect 3902 11526 3914 11586
rect 3914 11526 3964 11586
rect 3636 11524 3700 11526
rect 3724 11524 3788 11526
rect 3812 11524 3876 11526
rect 3900 11524 3964 11526
rect 10836 11586 10900 11588
rect 10924 11586 10988 11588
rect 11012 11586 11076 11588
rect 11100 11586 11164 11588
rect 10836 11526 10886 11586
rect 10886 11526 10898 11586
rect 10898 11526 10900 11586
rect 10924 11526 10958 11586
rect 10958 11526 10970 11586
rect 10970 11526 10988 11586
rect 11012 11526 11030 11586
rect 11030 11526 11042 11586
rect 11042 11526 11076 11586
rect 11100 11526 11102 11586
rect 11102 11526 11114 11586
rect 11114 11526 11164 11586
rect 10836 11524 10900 11526
rect 10924 11524 10988 11526
rect 11012 11524 11076 11526
rect 11100 11524 11164 11526
rect 18036 11586 18100 11588
rect 18124 11586 18188 11588
rect 18212 11586 18276 11588
rect 18300 11586 18364 11588
rect 18036 11526 18086 11586
rect 18086 11526 18098 11586
rect 18098 11526 18100 11586
rect 18124 11526 18158 11586
rect 18158 11526 18170 11586
rect 18170 11526 18188 11586
rect 18212 11526 18230 11586
rect 18230 11526 18242 11586
rect 18242 11526 18276 11586
rect 18300 11526 18302 11586
rect 18302 11526 18314 11586
rect 18314 11526 18364 11586
rect 18036 11524 18100 11526
rect 18124 11524 18188 11526
rect 18212 11524 18276 11526
rect 18300 11524 18364 11526
rect 25236 11586 25300 11588
rect 25324 11586 25388 11588
rect 25412 11586 25476 11588
rect 25500 11586 25564 11588
rect 25236 11526 25286 11586
rect 25286 11526 25298 11586
rect 25298 11526 25300 11586
rect 25324 11526 25358 11586
rect 25358 11526 25370 11586
rect 25370 11526 25388 11586
rect 25412 11526 25430 11586
rect 25430 11526 25442 11586
rect 25442 11526 25476 11586
rect 25500 11526 25502 11586
rect 25502 11526 25514 11586
rect 25514 11526 25564 11586
rect 25236 11524 25300 11526
rect 25324 11524 25388 11526
rect 25412 11524 25476 11526
rect 25500 11524 25564 11526
rect 32436 11585 32500 11587
rect 32524 11585 32588 11587
rect 32612 11585 32676 11587
rect 32700 11585 32764 11587
rect 32436 11525 32486 11585
rect 32486 11525 32498 11585
rect 32498 11525 32500 11585
rect 32524 11525 32558 11585
rect 32558 11525 32570 11585
rect 32570 11525 32588 11585
rect 32612 11525 32630 11585
rect 32630 11525 32642 11585
rect 32642 11525 32676 11585
rect 32700 11525 32702 11585
rect 32702 11525 32714 11585
rect 32714 11525 32764 11585
rect 32436 11523 32500 11525
rect 32524 11523 32588 11525
rect 32612 11523 32676 11525
rect 32700 11523 32764 11525
rect 3636 9410 3700 9412
rect 3724 9410 3788 9412
rect 3812 9410 3876 9412
rect 3900 9410 3964 9412
rect 3636 9350 3686 9410
rect 3686 9350 3698 9410
rect 3698 9350 3700 9410
rect 3724 9350 3758 9410
rect 3758 9350 3770 9410
rect 3770 9350 3788 9410
rect 3812 9350 3830 9410
rect 3830 9350 3842 9410
rect 3842 9350 3876 9410
rect 3900 9350 3902 9410
rect 3902 9350 3914 9410
rect 3914 9350 3964 9410
rect 3636 9348 3700 9350
rect 3724 9348 3788 9350
rect 3812 9348 3876 9350
rect 3900 9348 3964 9350
rect 10836 9410 10900 9412
rect 10924 9410 10988 9412
rect 11012 9410 11076 9412
rect 11100 9410 11164 9412
rect 10836 9350 10886 9410
rect 10886 9350 10898 9410
rect 10898 9350 10900 9410
rect 10924 9350 10958 9410
rect 10958 9350 10970 9410
rect 10970 9350 10988 9410
rect 11012 9350 11030 9410
rect 11030 9350 11042 9410
rect 11042 9350 11076 9410
rect 11100 9350 11102 9410
rect 11102 9350 11114 9410
rect 11114 9350 11164 9410
rect 10836 9348 10900 9350
rect 10924 9348 10988 9350
rect 11012 9348 11076 9350
rect 11100 9348 11164 9350
rect 18036 9410 18100 9412
rect 18124 9410 18188 9412
rect 18212 9410 18276 9412
rect 18300 9410 18364 9412
rect 18036 9350 18086 9410
rect 18086 9350 18098 9410
rect 18098 9350 18100 9410
rect 18124 9350 18158 9410
rect 18158 9350 18170 9410
rect 18170 9350 18188 9410
rect 18212 9350 18230 9410
rect 18230 9350 18242 9410
rect 18242 9350 18276 9410
rect 18300 9350 18302 9410
rect 18302 9350 18314 9410
rect 18314 9350 18364 9410
rect 18036 9348 18100 9350
rect 18124 9348 18188 9350
rect 18212 9348 18276 9350
rect 18300 9348 18364 9350
rect 25236 9410 25300 9412
rect 25324 9410 25388 9412
rect 25412 9410 25476 9412
rect 25500 9410 25564 9412
rect 25236 9350 25286 9410
rect 25286 9350 25298 9410
rect 25298 9350 25300 9410
rect 25324 9350 25358 9410
rect 25358 9350 25370 9410
rect 25370 9350 25388 9410
rect 25412 9350 25430 9410
rect 25430 9350 25442 9410
rect 25442 9350 25476 9410
rect 25500 9350 25502 9410
rect 25502 9350 25514 9410
rect 25514 9350 25564 9410
rect 25236 9348 25300 9350
rect 25324 9348 25388 9350
rect 25412 9348 25476 9350
rect 25500 9348 25564 9350
rect 32436 9410 32500 9412
rect 32524 9410 32588 9412
rect 32612 9410 32676 9412
rect 32700 9410 32764 9412
rect 32436 9350 32486 9410
rect 32486 9350 32498 9410
rect 32498 9350 32500 9410
rect 32524 9350 32558 9410
rect 32558 9350 32570 9410
rect 32570 9350 32588 9410
rect 32612 9350 32630 9410
rect 32630 9350 32642 9410
rect 32642 9350 32676 9410
rect 32700 9350 32702 9410
rect 32702 9350 32714 9410
rect 32714 9350 32764 9410
rect 32436 9348 32500 9350
rect 32524 9348 32588 9350
rect 32612 9348 32676 9350
rect 32700 9348 32764 9350
rect 3636 7234 3700 7236
rect 3724 7234 3788 7236
rect 3812 7234 3876 7236
rect 3900 7234 3964 7236
rect 3636 7174 3686 7234
rect 3686 7174 3698 7234
rect 3698 7174 3700 7234
rect 3724 7174 3758 7234
rect 3758 7174 3770 7234
rect 3770 7174 3788 7234
rect 3812 7174 3830 7234
rect 3830 7174 3842 7234
rect 3842 7174 3876 7234
rect 3900 7174 3902 7234
rect 3902 7174 3914 7234
rect 3914 7174 3964 7234
rect 3636 7172 3700 7174
rect 3724 7172 3788 7174
rect 3812 7172 3876 7174
rect 3900 7172 3964 7174
rect 10836 7234 10900 7236
rect 10924 7234 10988 7236
rect 11012 7234 11076 7236
rect 11100 7234 11164 7236
rect 10836 7174 10886 7234
rect 10886 7174 10898 7234
rect 10898 7174 10900 7234
rect 10924 7174 10958 7234
rect 10958 7174 10970 7234
rect 10970 7174 10988 7234
rect 11012 7174 11030 7234
rect 11030 7174 11042 7234
rect 11042 7174 11076 7234
rect 11100 7174 11102 7234
rect 11102 7174 11114 7234
rect 11114 7174 11164 7234
rect 10836 7172 10900 7174
rect 10924 7172 10988 7174
rect 11012 7172 11076 7174
rect 11100 7172 11164 7174
rect 25236 7234 25300 7236
rect 25324 7234 25388 7236
rect 25412 7234 25476 7236
rect 25500 7234 25564 7236
rect 25236 7174 25286 7234
rect 25286 7174 25298 7234
rect 25298 7174 25300 7234
rect 25324 7174 25358 7234
rect 25358 7174 25370 7234
rect 25370 7174 25388 7234
rect 25412 7174 25430 7234
rect 25430 7174 25442 7234
rect 25442 7174 25476 7234
rect 25500 7174 25502 7234
rect 25502 7174 25514 7234
rect 25514 7174 25564 7234
rect 25236 7172 25300 7174
rect 25324 7172 25388 7174
rect 25412 7172 25476 7174
rect 25500 7172 25564 7174
rect 32436 7234 32500 7236
rect 32524 7234 32588 7236
rect 32612 7234 32676 7236
rect 32700 7234 32764 7236
rect 32436 7174 32486 7234
rect 32486 7174 32498 7234
rect 32498 7174 32500 7234
rect 32524 7174 32558 7234
rect 32558 7174 32570 7234
rect 32570 7174 32588 7234
rect 32612 7174 32630 7234
rect 32630 7174 32642 7234
rect 32642 7174 32676 7234
rect 32700 7174 32702 7234
rect 32702 7174 32714 7234
rect 32714 7174 32764 7234
rect 32436 7172 32500 7174
rect 32524 7172 32588 7174
rect 32612 7172 32676 7174
rect 32700 7172 32764 7174
rect 7236 6280 7300 6282
rect 7324 6280 7388 6282
rect 7412 6280 7476 6282
rect 7500 6280 7564 6282
rect 7236 6220 7286 6280
rect 7286 6220 7298 6280
rect 7298 6220 7300 6280
rect 7324 6220 7358 6280
rect 7358 6220 7370 6280
rect 7370 6220 7388 6280
rect 7412 6220 7430 6280
rect 7430 6220 7442 6280
rect 7442 6220 7476 6280
rect 7500 6220 7502 6280
rect 7502 6220 7514 6280
rect 7514 6220 7564 6280
rect 7236 6218 7300 6220
rect 7324 6218 7388 6220
rect 7412 6218 7476 6220
rect 7500 6218 7564 6220
rect 14436 6280 14500 6282
rect 14524 6280 14588 6282
rect 14612 6280 14676 6282
rect 14700 6280 14764 6282
rect 14436 6220 14486 6280
rect 14486 6220 14498 6280
rect 14498 6220 14500 6280
rect 14524 6220 14558 6280
rect 14558 6220 14570 6280
rect 14570 6220 14588 6280
rect 14612 6220 14630 6280
rect 14630 6220 14642 6280
rect 14642 6220 14676 6280
rect 14700 6220 14702 6280
rect 14702 6220 14714 6280
rect 14714 6220 14764 6280
rect 14436 6218 14500 6220
rect 14524 6218 14588 6220
rect 14612 6218 14676 6220
rect 14700 6218 14764 6220
rect 21636 6280 21700 6282
rect 21724 6280 21788 6282
rect 21812 6280 21876 6282
rect 21900 6280 21964 6282
rect 21636 6220 21686 6280
rect 21686 6220 21698 6280
rect 21698 6220 21700 6280
rect 21724 6220 21758 6280
rect 21758 6220 21770 6280
rect 21770 6220 21788 6280
rect 21812 6220 21830 6280
rect 21830 6220 21842 6280
rect 21842 6220 21876 6280
rect 21900 6220 21902 6280
rect 21902 6220 21914 6280
rect 21914 6220 21964 6280
rect 21636 6218 21700 6220
rect 21724 6218 21788 6220
rect 21812 6218 21876 6220
rect 21900 6218 21964 6220
rect 28836 6280 28900 6282
rect 28924 6280 28988 6282
rect 29012 6280 29076 6282
rect 29100 6280 29164 6282
rect 28836 6220 28886 6280
rect 28886 6220 28898 6280
rect 28898 6220 28900 6280
rect 28924 6220 28958 6280
rect 28958 6220 28970 6280
rect 28970 6220 28988 6280
rect 29012 6220 29030 6280
rect 29030 6220 29042 6280
rect 29042 6220 29076 6280
rect 29100 6220 29102 6280
rect 29102 6220 29114 6280
rect 29114 6220 29164 6280
rect 28836 6218 28900 6220
rect 28924 6218 28988 6220
rect 29012 6218 29076 6220
rect 29100 6218 29164 6220
<< metal3 >>
rect 30602 20600 31602 21000
rect 30603 19800 31603 20200
rect 7200 14687 7600 14700
rect 7200 14614 7232 14687
rect 7304 14614 7320 14687
rect 7392 14614 7408 14687
rect 7480 14614 7496 14687
rect 7568 14614 7600 14687
rect 7200 14600 7600 14614
rect 14400 14687 14800 14700
rect 14400 14614 14432 14687
rect 14504 14614 14520 14687
rect 14592 14614 14608 14687
rect 14680 14614 14696 14687
rect 14768 14614 14800 14687
rect 14400 14600 14800 14614
rect 21600 14687 22000 14700
rect 21600 14614 21632 14687
rect 21704 14614 21720 14687
rect 21792 14614 21808 14687
rect 21880 14614 21896 14687
rect 21968 14614 22000 14687
rect 21600 14600 22000 14614
rect 28800 14687 29200 14700
rect 28800 14614 28832 14687
rect 28904 14614 28920 14687
rect 28992 14614 29008 14687
rect 29080 14614 29096 14687
rect 29168 14614 29200 14687
rect 28800 14600 29200 14614
rect 3600 13768 4000 13780
rect 3600 13696 3632 13768
rect 3704 13696 3720 13768
rect 3792 13696 3808 13768
rect 3880 13696 3896 13768
rect 3968 13696 4000 13768
rect 3600 13684 4000 13696
rect 10800 13768 11200 13780
rect 10800 13696 10832 13768
rect 10904 13696 10920 13768
rect 10992 13696 11008 13768
rect 11080 13696 11096 13768
rect 11168 13696 11200 13768
rect 10800 13684 11200 13696
rect 18000 13768 18400 13780
rect 18000 13696 18032 13768
rect 18104 13696 18120 13768
rect 18192 13696 18208 13768
rect 18280 13696 18296 13768
rect 18368 13696 18400 13768
rect 18000 13684 18400 13696
rect 25200 13768 25600 13780
rect 25200 13696 25232 13768
rect 25304 13696 25320 13768
rect 25392 13696 25408 13768
rect 25480 13696 25496 13768
rect 25568 13696 25600 13768
rect 25200 13684 25600 13696
rect 32400 13768 32800 13780
rect 32400 13696 32432 13768
rect 32504 13696 32520 13768
rect 32592 13696 32608 13768
rect 32680 13696 32696 13768
rect 32768 13696 32800 13768
rect 32400 13684 32800 13696
rect 3600 12680 4000 12692
rect 470 12420 542 12636
rect 3600 12608 3632 12680
rect 3704 12608 3720 12680
rect 3792 12608 3808 12680
rect 3880 12608 3896 12680
rect 3968 12608 4000 12680
rect 3600 12596 4000 12608
rect 470 12360 476 12420
rect 536 12360 542 12420
rect 470 12354 542 12360
rect 0 12137 400 12148
rect 0 12064 32 12137
rect 104 12064 120 12137
rect 192 12064 208 12137
rect 280 12064 296 12137
rect 368 12064 400 12137
rect 0 12052 400 12064
rect 36000 12137 36400 12148
rect 36000 12064 36032 12137
rect 36104 12064 36120 12137
rect 36192 12064 36208 12137
rect 36280 12064 36296 12137
rect 36368 12064 36400 12137
rect 36000 12052 36400 12064
rect 3600 11592 4000 11604
rect 3600 11520 3632 11592
rect 3704 11520 3720 11592
rect 3792 11520 3808 11592
rect 3880 11520 3896 11592
rect 3968 11520 4000 11592
rect 3600 11508 4000 11520
rect 10800 11592 11200 11604
rect 10800 11520 10832 11592
rect 10904 11520 10920 11592
rect 10992 11520 11008 11592
rect 11080 11520 11096 11592
rect 11168 11520 11200 11592
rect 10800 11508 11200 11520
rect 18000 11592 18400 11604
rect 18000 11520 18032 11592
rect 18104 11520 18120 11592
rect 18192 11520 18208 11592
rect 18280 11520 18296 11592
rect 18368 11520 18400 11592
rect 18000 11508 18400 11520
rect 25200 11592 25600 11604
rect 25200 11520 25232 11592
rect 25304 11520 25320 11592
rect 25392 11520 25408 11592
rect 25480 11520 25496 11592
rect 25568 11520 25600 11592
rect 25200 11508 25600 11520
rect 32400 11592 32800 11604
rect 32400 11519 32432 11592
rect 32504 11519 32520 11592
rect 32592 11519 32608 11592
rect 32680 11519 32696 11592
rect 32768 11519 32800 11592
rect 32400 11507 32800 11519
rect 3600 9417 4000 9428
rect 3600 9344 3632 9417
rect 3704 9344 3720 9417
rect 3792 9344 3808 9417
rect 3880 9344 3896 9417
rect 3968 9344 4000 9417
rect 3600 9332 4000 9344
rect 10800 9417 11200 9428
rect 10800 9344 10832 9417
rect 10904 9344 10920 9417
rect 10992 9344 11008 9417
rect 11080 9344 11096 9417
rect 11168 9344 11200 9417
rect 10800 9332 11200 9344
rect 18000 9417 18400 9428
rect 18000 9344 18032 9417
rect 18104 9344 18120 9417
rect 18192 9344 18208 9417
rect 18280 9344 18296 9417
rect 18368 9344 18400 9417
rect 18000 9332 18400 9344
rect 25200 9417 25600 9428
rect 25200 9344 25232 9417
rect 25304 9344 25320 9417
rect 25392 9344 25408 9417
rect 25480 9344 25496 9417
rect 25568 9344 25600 9417
rect 25200 9332 25600 9344
rect 32400 9417 32800 9428
rect 32400 9344 32432 9417
rect 32504 9344 32520 9417
rect 32592 9344 32608 9417
rect 32680 9344 32696 9417
rect 32768 9344 32800 9417
rect 32400 9332 32800 9344
rect 3600 7241 4000 7252
rect 3600 7168 3632 7241
rect 3704 7168 3720 7241
rect 3792 7168 3808 7241
rect 3880 7168 3896 7241
rect 3968 7168 4000 7241
rect 3600 7156 4000 7168
rect 10800 7241 11200 7252
rect 10800 7168 10832 7241
rect 10904 7168 10920 7241
rect 10992 7168 11008 7241
rect 11080 7168 11096 7241
rect 11168 7168 11200 7241
rect 10800 7156 11200 7168
rect 25200 7241 25600 7252
rect 25200 7168 25232 7241
rect 25304 7168 25320 7241
rect 25392 7168 25408 7241
rect 25480 7168 25496 7241
rect 25568 7168 25600 7241
rect 25200 7156 25600 7168
rect 32400 7241 32800 7252
rect 32400 7168 32432 7241
rect 32504 7168 32520 7241
rect 32592 7168 32608 7241
rect 32680 7168 32696 7241
rect 32768 7168 32800 7241
rect 32400 7156 32800 7168
rect 7200 6287 7600 6300
rect 7200 6214 7232 6287
rect 7304 6214 7320 6287
rect 7392 6214 7408 6287
rect 7480 6214 7496 6287
rect 7568 6214 7600 6287
rect 7200 6212 7600 6214
rect 14400 6287 14800 6300
rect 14400 6214 14432 6287
rect 14504 6214 14520 6287
rect 14592 6214 14608 6287
rect 14680 6214 14696 6287
rect 14768 6214 14800 6287
rect 7200 6200 7528 6212
rect 14400 6200 14800 6214
rect 21600 6287 22000 6300
rect 21600 6214 21632 6287
rect 21704 6214 21720 6287
rect 21792 6214 21808 6287
rect 21880 6214 21896 6287
rect 21968 6214 22000 6287
rect 21600 6200 22000 6214
rect 28800 6287 29200 6300
rect 28800 6214 28832 6287
rect 28904 6214 28920 6287
rect 28992 6214 29008 6287
rect 29080 6214 29096 6287
rect 29168 6214 29200 6287
rect 28800 6200 29200 6214
<< via3 >>
rect 7232 14682 7304 14687
rect 7232 14618 7236 14682
rect 7236 14618 7300 14682
rect 7300 14618 7304 14682
rect 7232 14614 7304 14618
rect 7320 14682 7392 14687
rect 7320 14618 7324 14682
rect 7324 14618 7388 14682
rect 7388 14618 7392 14682
rect 7320 14614 7392 14618
rect 7408 14682 7480 14687
rect 7408 14618 7412 14682
rect 7412 14618 7476 14682
rect 7476 14618 7480 14682
rect 7408 14614 7480 14618
rect 7496 14682 7568 14687
rect 7496 14618 7500 14682
rect 7500 14618 7564 14682
rect 7564 14618 7568 14682
rect 7496 14614 7568 14618
rect 14432 14682 14504 14687
rect 14432 14618 14436 14682
rect 14436 14618 14500 14682
rect 14500 14618 14504 14682
rect 14432 14614 14504 14618
rect 14520 14682 14592 14687
rect 14520 14618 14524 14682
rect 14524 14618 14588 14682
rect 14588 14618 14592 14682
rect 14520 14614 14592 14618
rect 14608 14682 14680 14687
rect 14608 14618 14612 14682
rect 14612 14618 14676 14682
rect 14676 14618 14680 14682
rect 14608 14614 14680 14618
rect 14696 14682 14768 14687
rect 14696 14618 14700 14682
rect 14700 14618 14764 14682
rect 14764 14618 14768 14682
rect 14696 14614 14768 14618
rect 21632 14682 21704 14687
rect 21632 14618 21636 14682
rect 21636 14618 21700 14682
rect 21700 14618 21704 14682
rect 21632 14614 21704 14618
rect 21720 14682 21792 14687
rect 21720 14618 21724 14682
rect 21724 14618 21788 14682
rect 21788 14618 21792 14682
rect 21720 14614 21792 14618
rect 21808 14682 21880 14687
rect 21808 14618 21812 14682
rect 21812 14618 21876 14682
rect 21876 14618 21880 14682
rect 21808 14614 21880 14618
rect 21896 14682 21968 14687
rect 21896 14618 21900 14682
rect 21900 14618 21964 14682
rect 21964 14618 21968 14682
rect 21896 14614 21968 14618
rect 28832 14682 28904 14687
rect 28832 14618 28836 14682
rect 28836 14618 28900 14682
rect 28900 14618 28904 14682
rect 28832 14614 28904 14618
rect 28920 14682 28992 14687
rect 28920 14618 28924 14682
rect 28924 14618 28988 14682
rect 28988 14618 28992 14682
rect 28920 14614 28992 14618
rect 29008 14682 29080 14687
rect 29008 14618 29012 14682
rect 29012 14618 29076 14682
rect 29076 14618 29080 14682
rect 29008 14614 29080 14618
rect 29096 14682 29168 14687
rect 29096 14618 29100 14682
rect 29100 14618 29164 14682
rect 29164 14618 29168 14682
rect 29096 14614 29168 14618
rect 3632 13764 3704 13768
rect 3632 13700 3636 13764
rect 3636 13700 3700 13764
rect 3700 13700 3704 13764
rect 3632 13696 3704 13700
rect 3720 13764 3792 13768
rect 3720 13700 3724 13764
rect 3724 13700 3788 13764
rect 3788 13700 3792 13764
rect 3720 13696 3792 13700
rect 3808 13764 3880 13768
rect 3808 13700 3812 13764
rect 3812 13700 3876 13764
rect 3876 13700 3880 13764
rect 3808 13696 3880 13700
rect 3896 13764 3968 13768
rect 3896 13700 3900 13764
rect 3900 13700 3964 13764
rect 3964 13700 3968 13764
rect 3896 13696 3968 13700
rect 10832 13764 10904 13768
rect 10832 13700 10836 13764
rect 10836 13700 10900 13764
rect 10900 13700 10904 13764
rect 10832 13696 10904 13700
rect 10920 13764 10992 13768
rect 10920 13700 10924 13764
rect 10924 13700 10988 13764
rect 10988 13700 10992 13764
rect 10920 13696 10992 13700
rect 11008 13764 11080 13768
rect 11008 13700 11012 13764
rect 11012 13700 11076 13764
rect 11076 13700 11080 13764
rect 11008 13696 11080 13700
rect 11096 13764 11168 13768
rect 11096 13700 11100 13764
rect 11100 13700 11164 13764
rect 11164 13700 11168 13764
rect 11096 13696 11168 13700
rect 18032 13764 18104 13768
rect 18032 13700 18036 13764
rect 18036 13700 18100 13764
rect 18100 13700 18104 13764
rect 18032 13696 18104 13700
rect 18120 13764 18192 13768
rect 18120 13700 18124 13764
rect 18124 13700 18188 13764
rect 18188 13700 18192 13764
rect 18120 13696 18192 13700
rect 18208 13764 18280 13768
rect 18208 13700 18212 13764
rect 18212 13700 18276 13764
rect 18276 13700 18280 13764
rect 18208 13696 18280 13700
rect 18296 13764 18368 13768
rect 18296 13700 18300 13764
rect 18300 13700 18364 13764
rect 18364 13700 18368 13764
rect 18296 13696 18368 13700
rect 25232 13764 25304 13768
rect 25232 13700 25236 13764
rect 25236 13700 25300 13764
rect 25300 13700 25304 13764
rect 25232 13696 25304 13700
rect 25320 13764 25392 13768
rect 25320 13700 25324 13764
rect 25324 13700 25388 13764
rect 25388 13700 25392 13764
rect 25320 13696 25392 13700
rect 25408 13764 25480 13768
rect 25408 13700 25412 13764
rect 25412 13700 25476 13764
rect 25476 13700 25480 13764
rect 25408 13696 25480 13700
rect 25496 13764 25568 13768
rect 25496 13700 25500 13764
rect 25500 13700 25564 13764
rect 25564 13700 25568 13764
rect 25496 13696 25568 13700
rect 32432 13764 32504 13768
rect 32432 13700 32436 13764
rect 32436 13700 32500 13764
rect 32500 13700 32504 13764
rect 32432 13696 32504 13700
rect 32520 13764 32592 13768
rect 32520 13700 32524 13764
rect 32524 13700 32588 13764
rect 32588 13700 32592 13764
rect 32520 13696 32592 13700
rect 32608 13764 32680 13768
rect 32608 13700 32612 13764
rect 32612 13700 32676 13764
rect 32676 13700 32680 13764
rect 32608 13696 32680 13700
rect 32696 13764 32768 13768
rect 32696 13700 32700 13764
rect 32700 13700 32764 13764
rect 32764 13700 32768 13764
rect 32696 13696 32768 13700
rect 3632 12676 3704 12680
rect 3632 12612 3636 12676
rect 3636 12612 3700 12676
rect 3700 12612 3704 12676
rect 3632 12608 3704 12612
rect 3720 12676 3792 12680
rect 3720 12612 3724 12676
rect 3724 12612 3788 12676
rect 3788 12612 3792 12676
rect 3720 12608 3792 12612
rect 3808 12676 3880 12680
rect 3808 12612 3812 12676
rect 3812 12612 3876 12676
rect 3876 12612 3880 12676
rect 3808 12608 3880 12612
rect 3896 12676 3968 12680
rect 3896 12612 3900 12676
rect 3900 12612 3964 12676
rect 3964 12612 3968 12676
rect 3896 12608 3968 12612
rect 32 12132 104 12137
rect 32 12068 36 12132
rect 36 12068 100 12132
rect 100 12068 104 12132
rect 32 12064 104 12068
rect 120 12132 192 12137
rect 120 12068 124 12132
rect 124 12068 188 12132
rect 188 12068 192 12132
rect 120 12064 192 12068
rect 208 12132 280 12137
rect 208 12068 212 12132
rect 212 12068 276 12132
rect 276 12068 280 12132
rect 208 12064 280 12068
rect 296 12132 368 12137
rect 296 12068 300 12132
rect 300 12068 364 12132
rect 364 12068 368 12132
rect 296 12064 368 12068
rect 36032 12132 36104 12137
rect 36032 12068 36036 12132
rect 36036 12068 36100 12132
rect 36100 12068 36104 12132
rect 36032 12064 36104 12068
rect 36120 12132 36192 12137
rect 36120 12068 36124 12132
rect 36124 12068 36188 12132
rect 36188 12068 36192 12132
rect 36120 12064 36192 12068
rect 36208 12132 36280 12137
rect 36208 12068 36212 12132
rect 36212 12068 36276 12132
rect 36276 12068 36280 12132
rect 36208 12064 36280 12068
rect 36296 12132 36368 12137
rect 36296 12068 36300 12132
rect 36300 12068 36364 12132
rect 36364 12068 36368 12132
rect 36296 12064 36368 12068
rect 3632 11588 3704 11592
rect 3632 11524 3636 11588
rect 3636 11524 3700 11588
rect 3700 11524 3704 11588
rect 3632 11520 3704 11524
rect 3720 11588 3792 11592
rect 3720 11524 3724 11588
rect 3724 11524 3788 11588
rect 3788 11524 3792 11588
rect 3720 11520 3792 11524
rect 3808 11588 3880 11592
rect 3808 11524 3812 11588
rect 3812 11524 3876 11588
rect 3876 11524 3880 11588
rect 3808 11520 3880 11524
rect 3896 11588 3968 11592
rect 3896 11524 3900 11588
rect 3900 11524 3964 11588
rect 3964 11524 3968 11588
rect 3896 11520 3968 11524
rect 10832 11588 10904 11592
rect 10832 11524 10836 11588
rect 10836 11524 10900 11588
rect 10900 11524 10904 11588
rect 10832 11520 10904 11524
rect 10920 11588 10992 11592
rect 10920 11524 10924 11588
rect 10924 11524 10988 11588
rect 10988 11524 10992 11588
rect 10920 11520 10992 11524
rect 11008 11588 11080 11592
rect 11008 11524 11012 11588
rect 11012 11524 11076 11588
rect 11076 11524 11080 11588
rect 11008 11520 11080 11524
rect 11096 11588 11168 11592
rect 11096 11524 11100 11588
rect 11100 11524 11164 11588
rect 11164 11524 11168 11588
rect 11096 11520 11168 11524
rect 18032 11588 18104 11592
rect 18032 11524 18036 11588
rect 18036 11524 18100 11588
rect 18100 11524 18104 11588
rect 18032 11520 18104 11524
rect 18120 11588 18192 11592
rect 18120 11524 18124 11588
rect 18124 11524 18188 11588
rect 18188 11524 18192 11588
rect 18120 11520 18192 11524
rect 18208 11588 18280 11592
rect 18208 11524 18212 11588
rect 18212 11524 18276 11588
rect 18276 11524 18280 11588
rect 18208 11520 18280 11524
rect 18296 11588 18368 11592
rect 18296 11524 18300 11588
rect 18300 11524 18364 11588
rect 18364 11524 18368 11588
rect 18296 11520 18368 11524
rect 25232 11588 25304 11592
rect 25232 11524 25236 11588
rect 25236 11524 25300 11588
rect 25300 11524 25304 11588
rect 25232 11520 25304 11524
rect 25320 11588 25392 11592
rect 25320 11524 25324 11588
rect 25324 11524 25388 11588
rect 25388 11524 25392 11588
rect 25320 11520 25392 11524
rect 25408 11588 25480 11592
rect 25408 11524 25412 11588
rect 25412 11524 25476 11588
rect 25476 11524 25480 11588
rect 25408 11520 25480 11524
rect 25496 11588 25568 11592
rect 25496 11524 25500 11588
rect 25500 11524 25564 11588
rect 25564 11524 25568 11588
rect 25496 11520 25568 11524
rect 32432 11587 32504 11592
rect 32432 11523 32436 11587
rect 32436 11523 32500 11587
rect 32500 11523 32504 11587
rect 32432 11519 32504 11523
rect 32520 11587 32592 11592
rect 32520 11523 32524 11587
rect 32524 11523 32588 11587
rect 32588 11523 32592 11587
rect 32520 11519 32592 11523
rect 32608 11587 32680 11592
rect 32608 11523 32612 11587
rect 32612 11523 32676 11587
rect 32676 11523 32680 11587
rect 32608 11519 32680 11523
rect 32696 11587 32768 11592
rect 32696 11523 32700 11587
rect 32700 11523 32764 11587
rect 32764 11523 32768 11587
rect 32696 11519 32768 11523
rect 3632 9412 3704 9417
rect 3632 9348 3636 9412
rect 3636 9348 3700 9412
rect 3700 9348 3704 9412
rect 3632 9344 3704 9348
rect 3720 9412 3792 9417
rect 3720 9348 3724 9412
rect 3724 9348 3788 9412
rect 3788 9348 3792 9412
rect 3720 9344 3792 9348
rect 3808 9412 3880 9417
rect 3808 9348 3812 9412
rect 3812 9348 3876 9412
rect 3876 9348 3880 9412
rect 3808 9344 3880 9348
rect 3896 9412 3968 9417
rect 3896 9348 3900 9412
rect 3900 9348 3964 9412
rect 3964 9348 3968 9412
rect 3896 9344 3968 9348
rect 10832 9412 10904 9417
rect 10832 9348 10836 9412
rect 10836 9348 10900 9412
rect 10900 9348 10904 9412
rect 10832 9344 10904 9348
rect 10920 9412 10992 9417
rect 10920 9348 10924 9412
rect 10924 9348 10988 9412
rect 10988 9348 10992 9412
rect 10920 9344 10992 9348
rect 11008 9412 11080 9417
rect 11008 9348 11012 9412
rect 11012 9348 11076 9412
rect 11076 9348 11080 9412
rect 11008 9344 11080 9348
rect 11096 9412 11168 9417
rect 11096 9348 11100 9412
rect 11100 9348 11164 9412
rect 11164 9348 11168 9412
rect 11096 9344 11168 9348
rect 18032 9412 18104 9417
rect 18032 9348 18036 9412
rect 18036 9348 18100 9412
rect 18100 9348 18104 9412
rect 18032 9344 18104 9348
rect 18120 9412 18192 9417
rect 18120 9348 18124 9412
rect 18124 9348 18188 9412
rect 18188 9348 18192 9412
rect 18120 9344 18192 9348
rect 18208 9412 18280 9417
rect 18208 9348 18212 9412
rect 18212 9348 18276 9412
rect 18276 9348 18280 9412
rect 18208 9344 18280 9348
rect 18296 9412 18368 9417
rect 18296 9348 18300 9412
rect 18300 9348 18364 9412
rect 18364 9348 18368 9412
rect 18296 9344 18368 9348
rect 25232 9412 25304 9417
rect 25232 9348 25236 9412
rect 25236 9348 25300 9412
rect 25300 9348 25304 9412
rect 25232 9344 25304 9348
rect 25320 9412 25392 9417
rect 25320 9348 25324 9412
rect 25324 9348 25388 9412
rect 25388 9348 25392 9412
rect 25320 9344 25392 9348
rect 25408 9412 25480 9417
rect 25408 9348 25412 9412
rect 25412 9348 25476 9412
rect 25476 9348 25480 9412
rect 25408 9344 25480 9348
rect 25496 9412 25568 9417
rect 25496 9348 25500 9412
rect 25500 9348 25564 9412
rect 25564 9348 25568 9412
rect 25496 9344 25568 9348
rect 32432 9412 32504 9417
rect 32432 9348 32436 9412
rect 32436 9348 32500 9412
rect 32500 9348 32504 9412
rect 32432 9344 32504 9348
rect 32520 9412 32592 9417
rect 32520 9348 32524 9412
rect 32524 9348 32588 9412
rect 32588 9348 32592 9412
rect 32520 9344 32592 9348
rect 32608 9412 32680 9417
rect 32608 9348 32612 9412
rect 32612 9348 32676 9412
rect 32676 9348 32680 9412
rect 32608 9344 32680 9348
rect 32696 9412 32768 9417
rect 32696 9348 32700 9412
rect 32700 9348 32764 9412
rect 32764 9348 32768 9412
rect 32696 9344 32768 9348
rect 3632 7236 3704 7241
rect 3632 7172 3636 7236
rect 3636 7172 3700 7236
rect 3700 7172 3704 7236
rect 3632 7168 3704 7172
rect 3720 7236 3792 7241
rect 3720 7172 3724 7236
rect 3724 7172 3788 7236
rect 3788 7172 3792 7236
rect 3720 7168 3792 7172
rect 3808 7236 3880 7241
rect 3808 7172 3812 7236
rect 3812 7172 3876 7236
rect 3876 7172 3880 7236
rect 3808 7168 3880 7172
rect 3896 7236 3968 7241
rect 3896 7172 3900 7236
rect 3900 7172 3964 7236
rect 3964 7172 3968 7236
rect 3896 7168 3968 7172
rect 10832 7236 10904 7241
rect 10832 7172 10836 7236
rect 10836 7172 10900 7236
rect 10900 7172 10904 7236
rect 10832 7168 10904 7172
rect 10920 7236 10992 7241
rect 10920 7172 10924 7236
rect 10924 7172 10988 7236
rect 10988 7172 10992 7236
rect 10920 7168 10992 7172
rect 11008 7236 11080 7241
rect 11008 7172 11012 7236
rect 11012 7172 11076 7236
rect 11076 7172 11080 7236
rect 11008 7168 11080 7172
rect 11096 7236 11168 7241
rect 11096 7172 11100 7236
rect 11100 7172 11164 7236
rect 11164 7172 11168 7236
rect 11096 7168 11168 7172
rect 25232 7236 25304 7241
rect 25232 7172 25236 7236
rect 25236 7172 25300 7236
rect 25300 7172 25304 7236
rect 25232 7168 25304 7172
rect 25320 7236 25392 7241
rect 25320 7172 25324 7236
rect 25324 7172 25388 7236
rect 25388 7172 25392 7236
rect 25320 7168 25392 7172
rect 25408 7236 25480 7241
rect 25408 7172 25412 7236
rect 25412 7172 25476 7236
rect 25476 7172 25480 7236
rect 25408 7168 25480 7172
rect 25496 7236 25568 7241
rect 25496 7172 25500 7236
rect 25500 7172 25564 7236
rect 25564 7172 25568 7236
rect 25496 7168 25568 7172
rect 32432 7236 32504 7241
rect 32432 7172 32436 7236
rect 32436 7172 32500 7236
rect 32500 7172 32504 7236
rect 32432 7168 32504 7172
rect 32520 7236 32592 7241
rect 32520 7172 32524 7236
rect 32524 7172 32588 7236
rect 32588 7172 32592 7236
rect 32520 7168 32592 7172
rect 32608 7236 32680 7241
rect 32608 7172 32612 7236
rect 32612 7172 32676 7236
rect 32676 7172 32680 7236
rect 32608 7168 32680 7172
rect 32696 7236 32768 7241
rect 32696 7172 32700 7236
rect 32700 7172 32764 7236
rect 32764 7172 32768 7236
rect 32696 7168 32768 7172
rect 7232 6282 7304 6287
rect 7232 6218 7236 6282
rect 7236 6218 7300 6282
rect 7300 6218 7304 6282
rect 7232 6214 7304 6218
rect 7320 6282 7392 6287
rect 7320 6218 7324 6282
rect 7324 6218 7388 6282
rect 7388 6218 7392 6282
rect 7320 6214 7392 6218
rect 7408 6282 7480 6287
rect 7408 6218 7412 6282
rect 7412 6218 7476 6282
rect 7476 6218 7480 6282
rect 7408 6214 7480 6218
rect 7496 6282 7568 6287
rect 7496 6218 7500 6282
rect 7500 6218 7564 6282
rect 7564 6218 7568 6282
rect 7496 6214 7568 6218
rect 14432 6282 14504 6287
rect 14432 6218 14436 6282
rect 14436 6218 14500 6282
rect 14500 6218 14504 6282
rect 14432 6214 14504 6218
rect 14520 6282 14592 6287
rect 14520 6218 14524 6282
rect 14524 6218 14588 6282
rect 14588 6218 14592 6282
rect 14520 6214 14592 6218
rect 14608 6282 14680 6287
rect 14608 6218 14612 6282
rect 14612 6218 14676 6282
rect 14676 6218 14680 6282
rect 14608 6214 14680 6218
rect 14696 6282 14768 6287
rect 14696 6218 14700 6282
rect 14700 6218 14764 6282
rect 14764 6218 14768 6282
rect 14696 6214 14768 6218
rect 21632 6282 21704 6287
rect 21632 6218 21636 6282
rect 21636 6218 21700 6282
rect 21700 6218 21704 6282
rect 21632 6214 21704 6218
rect 21720 6282 21792 6287
rect 21720 6218 21724 6282
rect 21724 6218 21788 6282
rect 21788 6218 21792 6282
rect 21720 6214 21792 6218
rect 21808 6282 21880 6287
rect 21808 6218 21812 6282
rect 21812 6218 21876 6282
rect 21876 6218 21880 6282
rect 21808 6214 21880 6218
rect 21896 6282 21968 6287
rect 21896 6218 21900 6282
rect 21900 6218 21964 6282
rect 21964 6218 21968 6282
rect 21896 6214 21968 6218
rect 28832 6282 28904 6287
rect 28832 6218 28836 6282
rect 28836 6218 28900 6282
rect 28900 6218 28904 6282
rect 28832 6214 28904 6218
rect 28920 6282 28992 6287
rect 28920 6218 28924 6282
rect 28924 6218 28988 6282
rect 28988 6218 28992 6282
rect 28920 6214 28992 6218
rect 29008 6282 29080 6287
rect 29008 6218 29012 6282
rect 29012 6218 29076 6282
rect 29076 6218 29080 6282
rect 29008 6214 29080 6218
rect 29096 6282 29168 6287
rect 29096 6218 29100 6282
rect 29100 6218 29164 6282
rect 29164 6218 29168 6282
rect 29096 6214 29168 6218
<< metal4 >>
rect 7200 14687 7600 14700
rect 7200 14614 7232 14687
rect 7304 14614 7320 14687
rect 7392 14614 7408 14687
rect 7480 14614 7496 14687
rect 7568 14614 7600 14687
rect 7200 14600 7600 14614
rect 14400 14687 14800 14700
rect 14400 14614 14432 14687
rect 14504 14614 14520 14687
rect 14592 14614 14608 14687
rect 14680 14614 14696 14687
rect 14768 14614 14800 14687
rect 14400 14600 14800 14614
rect 21600 14687 22000 14700
rect 21600 14614 21632 14687
rect 21704 14614 21720 14687
rect 21792 14614 21808 14687
rect 21880 14614 21896 14687
rect 21968 14614 22000 14687
rect 21600 14600 22000 14614
rect 28800 14687 29200 14700
rect 28800 14614 28832 14687
rect 28904 14614 28920 14687
rect 28992 14614 29008 14687
rect 29080 14614 29096 14687
rect 29168 14614 29200 14687
rect 28800 14600 29200 14614
rect 3600 13768 4000 13780
rect 3600 13696 3632 13768
rect 3704 13696 3720 13768
rect 3792 13696 3808 13768
rect 3880 13696 3896 13768
rect 3968 13696 4000 13768
rect 3600 13684 4000 13696
rect 10800 13768 11200 13780
rect 10800 13696 10832 13768
rect 10904 13696 10920 13768
rect 10992 13696 11008 13768
rect 11080 13696 11096 13768
rect 11168 13696 11200 13768
rect 10800 13684 11200 13696
rect 18000 13768 18400 13780
rect 18000 13696 18032 13768
rect 18104 13696 18120 13768
rect 18192 13696 18208 13768
rect 18280 13696 18296 13768
rect 18368 13696 18400 13768
rect 18000 13684 18400 13696
rect 25200 13768 25600 13780
rect 25200 13696 25232 13768
rect 25304 13696 25320 13768
rect 25392 13696 25408 13768
rect 25480 13696 25496 13768
rect 25568 13696 25600 13768
rect 25200 13684 25600 13696
rect 32400 13768 32800 13780
rect 32400 13696 32432 13768
rect 32504 13696 32520 13768
rect 32592 13696 32608 13768
rect 32680 13696 32696 13768
rect 32768 13696 32800 13768
rect 32400 13684 32800 13696
rect 3600 12680 4000 12692
rect 3600 12608 3632 12680
rect 3704 12608 3720 12680
rect 3792 12608 3808 12680
rect 3880 12608 3896 12680
rect 3968 12608 4000 12680
rect 3600 12596 4000 12608
rect 0 12137 400 12148
rect 0 12064 32 12137
rect 104 12064 120 12137
rect 192 12064 208 12137
rect 280 12064 296 12137
rect 368 12064 400 12137
rect 0 12052 400 12064
rect 36000 12137 36400 12148
rect 36000 12064 36032 12137
rect 36104 12064 36120 12137
rect 36192 12064 36208 12137
rect 36280 12064 36296 12137
rect 36368 12064 36400 12137
rect 36000 12052 36400 12064
rect 3600 11592 4000 11604
rect 3600 11520 3632 11592
rect 3704 11520 3720 11592
rect 3792 11520 3808 11592
rect 3880 11520 3896 11592
rect 3968 11520 4000 11592
rect 3600 11508 4000 11520
rect 10800 11592 11200 11604
rect 10800 11520 10832 11592
rect 10904 11520 10920 11592
rect 10992 11520 11008 11592
rect 11080 11520 11096 11592
rect 11168 11520 11200 11592
rect 10800 11508 11200 11520
rect 18000 11592 18400 11604
rect 18000 11520 18032 11592
rect 18104 11520 18120 11592
rect 18192 11520 18208 11592
rect 18280 11520 18296 11592
rect 18368 11520 18400 11592
rect 18000 11508 18400 11520
rect 25200 11592 25600 11604
rect 25200 11520 25232 11592
rect 25304 11520 25320 11592
rect 25392 11520 25408 11592
rect 25480 11520 25496 11592
rect 25568 11520 25600 11592
rect 25200 11508 25600 11520
rect 32400 11592 32800 11604
rect 32400 11519 32432 11592
rect 32504 11519 32520 11592
rect 32592 11519 32608 11592
rect 32680 11519 32696 11592
rect 32768 11519 32800 11592
rect 32400 11507 32800 11519
rect 3600 9417 4000 9428
rect 3600 9344 3632 9417
rect 3704 9344 3720 9417
rect 3792 9344 3808 9417
rect 3880 9344 3896 9417
rect 3968 9344 4000 9417
rect 3600 9332 4000 9344
rect 10800 9417 11200 9428
rect 10800 9344 10832 9417
rect 10904 9344 10920 9417
rect 10992 9344 11008 9417
rect 11080 9344 11096 9417
rect 11168 9344 11200 9417
rect 10800 9332 11200 9344
rect 18000 9417 18400 9428
rect 18000 9344 18032 9417
rect 18104 9344 18120 9417
rect 18192 9344 18208 9417
rect 18280 9344 18296 9417
rect 18368 9344 18400 9417
rect 18000 9332 18400 9344
rect 25200 9417 25600 9428
rect 25200 9344 25232 9417
rect 25304 9344 25320 9417
rect 25392 9344 25408 9417
rect 25480 9344 25496 9417
rect 25568 9344 25600 9417
rect 25200 9332 25600 9344
rect 32400 9417 32800 9428
rect 32400 9344 32432 9417
rect 32504 9344 32520 9417
rect 32592 9344 32608 9417
rect 32680 9344 32696 9417
rect 32768 9344 32800 9417
rect 32400 9332 32800 9344
rect 3600 7241 4000 7252
rect 3600 7168 3632 7241
rect 3704 7168 3720 7241
rect 3792 7168 3808 7241
rect 3880 7168 3896 7241
rect 3968 7168 4000 7241
rect 3600 7156 4000 7168
rect 10800 7241 11200 7252
rect 10800 7168 10832 7241
rect 10904 7168 10920 7241
rect 10992 7168 11008 7241
rect 11080 7168 11096 7241
rect 11168 7168 11200 7241
rect 10800 7156 11200 7168
rect 25200 7241 25600 7252
rect 25200 7168 25232 7241
rect 25304 7168 25320 7241
rect 25392 7168 25408 7241
rect 25480 7168 25496 7241
rect 25568 7168 25600 7241
rect 25200 7156 25600 7168
rect 32400 7241 32800 7252
rect 32400 7168 32432 7241
rect 32504 7168 32520 7241
rect 32592 7168 32608 7241
rect 32680 7168 32696 7241
rect 32768 7168 32800 7241
rect 32400 7156 32800 7168
rect 7200 6287 7600 6300
rect 7200 6214 7232 6287
rect 7304 6214 7320 6287
rect 7392 6214 7408 6287
rect 7480 6214 7496 6287
rect 7568 6214 7600 6287
rect 7200 6212 7600 6214
rect 14400 6287 14800 6300
rect 14400 6214 14432 6287
rect 14504 6214 14520 6287
rect 14592 6214 14608 6287
rect 14680 6214 14696 6287
rect 14768 6214 14800 6287
rect 7200 6200 7528 6212
rect 14400 6200 14800 6214
rect 21600 6287 22000 6300
rect 21600 6214 21632 6287
rect 21704 6214 21720 6287
rect 21792 6214 21808 6287
rect 21880 6214 21896 6287
rect 21968 6214 22000 6287
rect 21600 6200 22000 6214
rect 28800 6287 29200 6300
rect 28800 6214 28832 6287
rect 28904 6214 28920 6287
rect 28992 6214 29008 6287
rect 29080 6214 29096 6287
rect 29168 6214 29200 6287
rect 28800 6200 29200 6214
use ring_osc_r100  ring_osc_r100_0
timestamp 1624957116
transform 1 0 -98 0 1 6660
box 100 -58 36300 7674
use power_ring_2_2  power_ring_2_2_0
timestamp 1624938805
transform 1 0 -27000 0 1 -3200
box 27000 3200 63400 24200
use pwell_co_ring  pwell_co_ring_0
timestamp 1624938805
transform 1 0 -98 0 1 200
box 176 6000 36124 14500
<< labels >>
flabel locali 1229 12475 1398 12535 1 FreeSans 400 0 0 0 hi_logic
flabel metal1 30904 10962 31422 11060 1 FreeSans 2 0 0 0 v_crt
flabel metal1 9238 12852 9536 12980 1 FreeSans 2 0 0 0 pn[6]
flabel metal1 15150 12854 15448 12982 1 FreeSans 2 0 0 0 pn[7]
flabel metal1 21054 12852 21352 12980 1 FreeSans 2 0 0 0 pn[8]
flabel metal1 26946 12852 27244 12980 1 FreeSans 2 0 0 0 pn[9]
flabel metal1 29670 7954 29968 8082 1 FreeSans 2 0 0 0 pn[0]
flabel metal1 23754 7954 24052 8082 1 FreeSans 2 0 0 0 pn[1]
flabel metal1 17858 7954 18156 8082 1 FreeSans 2 0 0 0 pn[2]
flabel metal1 11946 7954 12244 8082 1 FreeSans 2 0 0 0 pn[3]
flabel metal1 6046 7956 6344 8084 1 FreeSans 2 0 0 0 pn[4]
flabel metal2 702 10532 1018 10670 1 FreeSans 2 0 0 0 pn[5]
flabel metal2 34266 10048 34582 10186 1 FreeSans 2 0 0 0 pn[10]
flabel locali 1688 12416 1732 12460 1 FreeSans 2 0 0 0 lo_logic
flabel metal2 36502 11738 36702 11898 1 FreeSans 2400 0 0 0 input_analog
port 12 nsew signal input
flabel metal3 s 30603 19800 31603 20200 1 FreeSans 2400 0 0 0 vssd2
port 14 nsew ground bidirectional abutment
flabel metal3 s 30602 20600 31602 21000 1 FreeSans 2400 0 0 0 vccd2
port 13 nsew power bidirectional abutment
flabel metal2 1228 8510 1412 8602 1 FreeSans 2000 0 0 0 p[0]
port 1 nsew signal output
flabel metal2 6118 8510 6302 8602 1 FreeSans 2000 0 0 0 p[1]
port 2 nsew signal output
flabel metal2 12006 8510 12190 8602 1 FreeSans 2000 0 0 0 p[3]
port 4 nsew signal output
flabel metal2 17894 8510 18078 8602 1 FreeSans 2000 0 0 0 p[5]
port 6 nsew signal output
flabel metal2 23874 8510 24058 8602 1 FreeSans 2000 0 0 0 p[7]
port 8 nsew signal output
flabel metal2 29762 8510 29946 8602 1 FreeSans 2000 0 0 0 p[9]
port 10 nsew signal output
flabel metal2 33166 8510 33350 8602 1 FreeSans 2000 0 0 0 p[10]
port 11 nsew signal output
flabel metal2 9246 12326 9430 12418 1 FreeSans 2000 0 0 0 p[2]
port 3 nsew signal output
flabel metal2 15134 12326 15318 12418 1 FreeSans 2000 0 0 0 p[4]
port 5 nsew signal output
flabel metal2 21022 12326 21206 12418 1 FreeSans 2000 0 0 0 p[6]
port 7 nsew signal output
flabel metal2 26910 12326 27094 12418 1 FreeSans 2000 0 0 0 p[8]
port 9 nsew signal output
flabel metal3 474 12438 534 12622 3 FreeSans 1600 90 0 0 enb
port 15 nsew signal input
<< end >>
