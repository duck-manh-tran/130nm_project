magic
tech sky130A
magscale 1 2
timestamp 1624688222
<< ndiff >>
rect 1627 12258 1661 12292
<< pdiff >>
rect 1627 12582 1661 12616
<< locali >>
rect 1910 12548 1955 12592
rect 2308 12542 2353 12586
rect 62 12438 158 12460
rect 62 12382 74 12438
rect 130 12406 158 12438
rect 130 12382 142 12406
rect 1496 12384 1521 12418
rect 62 12360 142 12382
<< viali >>
rect 74 12382 130 12438
<< metal1 >>
rect 0 12656 1994 12752
rect 62 12438 142 12484
rect 62 12382 74 12438
rect 130 12382 142 12438
rect 10568 12390 10574 12462
rect 10646 12390 10652 12462
rect 14110 12390 14116 12462
rect 14188 12390 14194 12462
rect 16656 12390 16662 12462
rect 16734 12390 16740 12462
rect 21082 12390 21170 12462
rect 21242 12390 21382 12462
rect 21722 12404 23600 12476
rect 62 12348 142 12382
rect 800 12112 1962 12208
rect 1226 8706 1390 8778
rect 1462 8706 1562 8778
rect 4774 8706 4780 8778
rect 4852 8706 4858 8778
rect 8560 8706 8566 8778
rect 8638 8706 8644 8778
rect 13160 8706 13166 8778
rect 13238 8706 13244 8778
rect 15644 8706 15650 8778
rect 15722 8706 15728 8778
rect 19232 8706 19238 8778
rect 19310 8706 19316 8778
<< via1 >>
rect 5898 12390 5970 12462
rect 10574 12390 10646 12462
rect 14116 12390 14188 12462
rect 16662 12390 16734 12462
rect 21170 12390 21242 12462
rect 1390 8706 1462 8778
rect 4780 8706 4852 8778
rect 8566 8706 8638 8778
rect 13166 8706 13238 8778
rect 15650 8706 15722 8778
rect 19238 8706 19310 8778
<< metal2 >>
rect 5842 12462 6026 12472
rect 5842 12390 5898 12462
rect 5970 12390 6026 12462
rect 5842 12380 6026 12390
rect 10518 12462 10702 12472
rect 10518 12390 10574 12462
rect 10646 12390 10702 12462
rect 10518 12380 10702 12390
rect 14060 12462 14244 12472
rect 14060 12390 14116 12462
rect 14188 12390 14244 12462
rect 14060 12380 14244 12390
rect 16606 12462 16790 12472
rect 16606 12390 16662 12462
rect 16734 12390 16790 12462
rect 16606 12380 16790 12390
rect 21114 12462 21298 12472
rect 21114 12390 21170 12462
rect 21242 12390 21298 12462
rect 21114 12380 21298 12390
rect 24426 11522 24610 11542
rect 24426 11462 24488 11522
rect 24548 11462 24610 11522
rect 24426 11442 24610 11462
rect 1334 8778 1518 8788
rect 1334 8706 1390 8778
rect 1462 8706 1518 8778
rect 1334 8696 1518 8706
rect 4724 8778 4908 8788
rect 4724 8706 4780 8778
rect 4852 8706 4908 8778
rect 4724 8696 4908 8706
rect 8510 8778 8694 8788
rect 8510 8706 8566 8778
rect 8638 8706 8694 8778
rect 8510 8696 8694 8706
rect 13110 8778 13294 8788
rect 13110 8706 13166 8778
rect 13238 8706 13294 8778
rect 13110 8696 13294 8706
rect 15594 8778 15778 8788
rect 15594 8706 15650 8778
rect 15722 8706 15778 8778
rect 15594 8696 15778 8706
rect 19182 8778 19366 8788
rect 19182 8706 19238 8778
rect 19310 8706 19366 8778
rect 19182 8696 19366 8706
<< via2 >>
rect 24488 11462 24548 11522
<< metal3 >>
rect 0 20600 5200 21000
rect 24464 11522 24572 11628
rect 24464 11462 24488 11522
rect 24548 11462 24572 11522
rect 24464 11356 24572 11462
rect 18600 800 23600 1200
use ring_osc_w6  ring_osc_w6_0
timestamp 1624684182
transform 1 0 1500 0 1 7600
box -1410 0 23110 5968
use via_m1  via_m1_4
timestamp 1623561200
transform 1 0 -7298 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_5
timestamp 1623561200
transform 1 0 -1698 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_8
timestamp 1623561200
transform 1 0 3902 0 1 662
box 10898 6956 11298 7052
use via_m1  via_m1_9
timestamp 1623561200
transform 1 0 9502 0 1 662
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_4
timestamp 1623563441
transform 1 0 6400 0 1 7360
box 0 2 400 98
use via_m4_li  via_m4_li_5
timestamp 1623563441
transform 1 0 12000 0 1 7360
box 0 2 400 98
use pwell_co_ring_w6  pwell_co_ring_w6_0
timestamp 1623529308
transform 1 0 3020 0 1 13740
box -1680 -6360 20145 60
use via_m1  via_m1_1
timestamp 1623561200
transform 1 0 -10898 0 1 5700
box 10898 6956 11298 7052
use via_m1  via_m1_2
timestamp 1623561200
transform 1 0 -10098 0 1 5156
box 10898 6956 11298 7052
use via_m1  via_m1_3
timestamp 1623561200
transform 1 0 -7298 0 1 6498
box 10898 6956 11298 7052
use via_m1  via_m1_6
timestamp 1623561200
transform 1 0 -1698 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_3
timestamp 1623563441
transform 1 0 6400 0 1 13720
box 0 2 400 98
use via_m1  via_m1_7
timestamp 1623561200
transform 1 0 3902 0 1 6498
box 10898 6956 11298 7052
use via_m4_li  via_m4_li_2
timestamp 1623563441
transform 1 0 12000 0 1 13720
box 0 2 400 98
use via_m4_li  via_m4_li_1
timestamp 1623563441
transform 1 0 17600 0 1 13720
box 0 2 400 98
use via_m1  via_m1_11
timestamp 1623561200
transform 1 0 12302 0 1 5436
box 10898 6956 11298 7052
use via_m1  via_m1_10
timestamp 1623561200
transform 1 0 9502 0 1 6498
box 10898 6956 11298 7052
use power_ring  power_ring_0
timestamp 1623530672
transform 1 0 0 0 1 0
box 0 0 24400 21000
<< labels >>
flabel metal3 0 20600 5200 21000 1 FreeSans 16 0 0 0 vccd2
port 14 n power bidirectional
flabel metal3 18600 800 23600 1200 1 FreeSans 16 0 0 0 vssd2
port 15 s ground bidirectional
flabel metal2 24468 11442 24568 11542 1 FreeSans 640 0 0 0 input_analog
port 13 e signal input
flabel metal1 62 12378 142 12458 1 FreeSans 640 0 0 0 enb
port 12 w signal input
flabel metal2 1384 8700 1468 8784 1 FreeSans 640 0 0 0 p[0]
port 6 s signal output
flabel metal2 8560 8700 8644 8784 1 FreeSans 640 0 0 0 p[3]
port 4 s signal output
flabel metal2 13160 8700 13244 8784 1 FreeSans 640 0 0 0 p[5]
port 3 s signal output
flabel metal2 15644 8700 15728 8784 1 FreeSans 640 0 0 0 p[7]
port 2 s signal output
flabel metal2 19232 8700 19316 8784 1 FreeSans 640 0 0 0 p[9]
port 1 s signal output
flabel metal2 14110 12384 14194 12468 1 FreeSans 640 0 0 0 p[6]
port 9 n signal output
flabel metal2 16656 12384 16740 12468 1 FreeSans 640 0 0 0 p[8]
port 10 nsew default output
flabel metal2 21164 12384 21248 12468 1 FreeSans 640 0 0 0 p[10]
port 11 n signal output
flabel metal2 4774 8700 4858 8784 1 FreeSans 640 0 0 0 p[1]
port 5 s signal output
flabel metal2 5892 12384 5976 12468 1 FreeSans 640 0 0 0 p[2]
port 7 n signal output
flabel metal2 10568 12384 10652 12468 1 FreeSans 640 0 0 0 p[4]
port 8 n signal output
<< end >>
50 41 62 33 74 25 86 17 98 0 10
