magic
tech sky130A
magscale 1 2
timestamp 1623172293
<< nwell >>
rect 726 6022 1262 6068
rect 1560 6022 1912 6068
rect 868 5998 1062 6022
rect 1668 5998 1862 6022
<< nsubdiff >>
rect 868 5998 904 6032
rect 944 5998 984 6032
rect 1024 5998 1062 6032
rect 1668 5998 1704 6032
rect 1744 5998 1784 6032
rect 1824 5998 1862 6032
<< nsubdiffcont >>
rect 904 5998 944 6032
rect 984 5998 1024 6032
rect 1704 5998 1744 6032
rect 1784 5998 1824 6032
<< locali >>
rect 868 5998 904 6032
rect 944 5998 984 6032
rect 1024 5998 1062 6032
rect 1668 5998 1704 6032
rect 1744 5998 1784 6032
rect 1824 5998 1862 6032
rect 1266 5831 1556 5875
rect 1159 5815 1556 5831
rect 1159 5771 1326 5815
rect 1496 5788 1556 5815
rect 1372 5729 1432 5742
rect 1372 5695 1385 5729
rect 1419 5695 1432 5729
rect 1496 5728 1663 5788
rect 807 5652 857 5685
rect 1372 5575 1432 5695
rect 1206 5515 1432 5575
<< viali >>
rect 1385 5695 1419 5729
<< metal1 >>
rect 3256 7568 3578 7664
rect 7800 7640 8000 7664
rect 7852 7588 7874 7640
rect 7926 7588 7948 7640
rect 7800 7568 8000 7588
rect 14000 7640 14200 7664
rect 14052 7588 14074 7640
rect 14126 7588 14148 7640
rect 14000 7568 14200 7588
rect 22400 7640 22600 7664
rect 22452 7588 22474 7640
rect 22526 7588 22548 7640
rect 22400 7568 22600 7588
rect 28600 7640 28800 7664
rect 28652 7588 28674 7640
rect 28726 7588 28748 7640
rect 28600 7568 28800 7588
rect 33078 7642 34698 7664
rect 33078 7590 34498 7642
rect 34550 7590 34562 7642
rect 34614 7590 34626 7642
rect 34678 7590 34698 7642
rect 33078 7568 34698 7590
rect 3200 7024 6778 7120
rect 3568 6315 3767 6323
rect 3568 6199 3609 6315
rect 3725 6199 3767 6315
rect 3568 6191 3767 6199
rect 9336 6192 9634 6320
rect 15248 6194 15546 6322
rect 21152 6192 21450 6320
rect 27044 6192 27342 6320
rect 32884 6315 33088 6323
rect 32884 6199 32896 6315
rect 33076 6199 33088 6315
rect 32884 6191 33088 6199
rect 1006 5936 4058 6032
rect 3400 5770 3783 5772
rect 1360 5742 1444 5748
rect 3400 5742 3585 5770
rect 1360 5729 3585 5742
rect 1360 5695 1385 5729
rect 1419 5695 3585 5729
rect 1360 5682 3585 5695
rect 1360 5676 1444 5682
rect 3400 5654 3585 5682
rect 3765 5654 3783 5770
rect 3400 5652 3783 5654
rect 9310 5770 9430 5772
rect 9310 5654 9312 5770
rect 9428 5654 9430 5770
rect 9310 5652 9430 5654
rect 9458 5770 9578 5772
rect 9458 5654 9460 5770
rect 9576 5654 9578 5770
rect 9458 5652 9578 5654
rect 15210 5770 15330 5772
rect 15210 5654 15212 5770
rect 15328 5654 15330 5770
rect 15210 5652 15330 5654
rect 15358 5770 15478 5772
rect 15358 5654 15360 5770
rect 15476 5654 15478 5770
rect 15358 5652 15478 5654
rect 21110 5770 21230 5772
rect 21110 5654 21112 5770
rect 21228 5654 21230 5770
rect 21110 5652 21230 5654
rect 21258 5770 21378 5772
rect 21258 5654 21260 5770
rect 21376 5654 21378 5770
rect 21258 5652 21378 5654
rect 27010 5770 27130 5772
rect 27010 5654 27012 5770
rect 27128 5654 27130 5770
rect 27010 5652 27130 5654
rect 27158 5770 27278 5772
rect 27158 5654 27160 5770
rect 27276 5654 27278 5770
rect 27158 5652 27278 5654
rect 32880 5770 33088 5772
rect 32880 5654 32894 5770
rect 33074 5654 33088 5770
rect 32880 5652 33088 5654
rect 0 5392 1993 5488
rect 3001 4848 6579 4944
rect 33078 4848 34488 4944
rect 7800 4398 8000 4400
rect 14000 4398 14200 4400
rect 22400 4398 22600 4400
rect 30842 4398 31260 4400
rect 3400 4382 35506 4398
rect 3400 4376 34631 4382
rect 3400 4324 7800 4376
rect 7852 4324 7874 4376
rect 7926 4324 7948 4376
rect 8000 4324 14000 4376
rect 14052 4324 14074 4376
rect 14126 4324 14148 4376
rect 14200 4324 22400 4376
rect 22452 4324 22474 4376
rect 22526 4324 22548 4376
rect 22600 4324 28600 4376
rect 28652 4324 28674 4376
rect 28726 4324 28748 4376
rect 28800 4330 34631 4376
rect 34683 4330 34706 4382
rect 34758 4330 34782 4382
rect 34834 4330 34857 4382
rect 34909 4330 34932 4382
rect 34984 4330 35007 4382
rect 35059 4330 35083 4382
rect 35135 4330 35158 4382
rect 35210 4330 35233 4382
rect 35285 4330 35307 4382
rect 35359 4330 35383 4382
rect 35435 4330 35506 4382
rect 28800 4324 35506 4330
rect 3400 4302 35506 4324
rect 7800 3288 8000 3312
rect 7852 3236 7874 3288
rect 7926 3236 7948 3288
rect 7800 3216 8000 3236
rect 14000 3288 14200 3312
rect 14052 3236 14074 3288
rect 14126 3236 14148 3288
rect 14000 3216 14200 3236
rect 22400 3288 22600 3312
rect 22452 3236 22474 3288
rect 22526 3236 22548 3288
rect 22400 3216 22600 3236
rect 28600 3288 28800 3312
rect 28652 3236 28674 3288
rect 28726 3236 28748 3288
rect 28600 3216 28800 3236
rect 35353 3290 36088 3312
rect 35353 3238 35893 3290
rect 35945 3238 35957 3290
rect 36009 3238 36021 3290
rect 36073 3238 36088 3290
rect 35353 3216 36088 3238
rect 0 2672 400 2768
rect 35353 2672 35888 2768
rect 1341 1962 1481 1964
rect 1341 1846 1353 1962
rect 1469 1846 1481 1962
rect 1341 1844 1481 1846
rect 6200 1962 6320 1964
rect 6200 1846 6202 1962
rect 6318 1846 6320 1962
rect 6200 1844 6320 1846
rect 6348 1962 6468 1964
rect 6348 1846 6350 1962
rect 6466 1846 6468 1962
rect 6348 1844 6468 1846
rect 12100 1962 12220 1964
rect 12100 1846 12102 1962
rect 12218 1846 12220 1962
rect 12100 1844 12220 1846
rect 12248 1962 12368 1964
rect 12248 1846 12250 1962
rect 12366 1846 12368 1962
rect 12248 1844 12368 1846
rect 18000 1962 18120 1964
rect 18000 1846 18002 1962
rect 18118 1846 18120 1962
rect 18000 1844 18120 1846
rect 18148 1962 18268 1964
rect 18148 1846 18150 1962
rect 18266 1846 18268 1962
rect 18148 1844 18268 1846
rect 23900 1962 24020 1964
rect 23900 1846 23902 1962
rect 24018 1846 24020 1962
rect 23900 1844 24020 1846
rect 24048 1962 24168 1964
rect 24048 1846 24050 1962
rect 24166 1846 24168 1962
rect 24048 1844 24168 1846
rect 29800 1962 29920 1964
rect 29800 1846 29802 1962
rect 29918 1846 29920 1962
rect 29800 1844 29920 1846
rect 29932 1962 30068 1964
rect 29932 1846 29950 1962
rect 30066 1846 30068 1962
rect 29932 1844 30068 1846
rect 33208 1962 33492 1964
rect 33208 1846 33230 1962
rect 33346 1846 33374 1962
rect 33490 1846 33492 1962
rect 33208 1844 33492 1846
rect 406 1294 704 1422
rect 789 1417 949 1425
rect 789 1301 811 1417
rect 927 1301 949 1417
rect 789 1293 949 1301
rect 6014 1293 6983 1425
rect 11914 1293 12883 1425
rect 17814 1293 18783 1425
rect 23714 1293 24683 1425
rect 29614 1293 30583 1425
rect 34528 1417 35366 1419
rect 34528 1301 34552 1417
rect 34668 1301 35366 1417
rect 34528 1299 35366 1301
rect 35502 1294 35800 1422
rect 0 496 400 592
rect 35353 496 35888 592
rect 7800 24 8000 48
rect 7852 -28 7874 24
rect 7926 -28 7948 24
rect 7800 -48 8000 -28
rect 14000 24 14200 48
rect 14052 -28 14074 24
rect 14126 -28 14148 24
rect 14000 -48 14200 -28
rect 22400 24 22600 48
rect 22452 -28 22474 24
rect 22526 -28 22548 24
rect 22400 -48 22600 -28
rect 28600 24 28800 48
rect 28652 -28 28674 24
rect 28726 -28 28748 24
rect 28600 -48 28800 -28
rect 35353 26 36088 48
rect 35353 -26 35895 26
rect 35947 -26 35959 26
rect 36011 -26 36023 26
rect 36075 -26 36088 26
rect 35353 -48 36088 -26
<< via1 >>
rect 7800 7588 7852 7640
rect 7874 7588 7926 7640
rect 7948 7588 8000 7640
rect 14000 7588 14052 7640
rect 14074 7588 14126 7640
rect 14148 7588 14200 7640
rect 22400 7588 22452 7640
rect 22474 7588 22526 7640
rect 22548 7588 22600 7640
rect 28600 7588 28652 7640
rect 28674 7588 28726 7640
rect 28748 7588 28800 7640
rect 34498 7590 34550 7642
rect 34562 7590 34614 7642
rect 34626 7590 34678 7642
rect 3609 6199 3725 6315
rect 32896 6199 33076 6315
rect 3585 5654 3765 5770
rect 9312 5654 9428 5770
rect 9460 5654 9576 5770
rect 15212 5654 15328 5770
rect 15360 5654 15476 5770
rect 21112 5654 21228 5770
rect 21260 5654 21376 5770
rect 27012 5654 27128 5770
rect 27160 5654 27276 5770
rect 32894 5654 33074 5770
rect 7800 4324 7852 4376
rect 7874 4324 7926 4376
rect 7948 4324 8000 4376
rect 14000 4324 14052 4376
rect 14074 4324 14126 4376
rect 14148 4324 14200 4376
rect 22400 4324 22452 4376
rect 22474 4324 22526 4376
rect 22548 4324 22600 4376
rect 28600 4324 28652 4376
rect 28674 4324 28726 4376
rect 28748 4324 28800 4376
rect 34631 4330 34683 4382
rect 34706 4330 34758 4382
rect 34782 4330 34834 4382
rect 34857 4330 34909 4382
rect 34932 4330 34984 4382
rect 35007 4330 35059 4382
rect 35083 4330 35135 4382
rect 35158 4330 35210 4382
rect 35233 4330 35285 4382
rect 35307 4330 35359 4382
rect 35383 4330 35435 4382
rect 7800 3236 7852 3288
rect 7874 3236 7926 3288
rect 7948 3236 8000 3288
rect 14000 3236 14052 3288
rect 14074 3236 14126 3288
rect 14148 3236 14200 3288
rect 22400 3236 22452 3288
rect 22474 3236 22526 3288
rect 22548 3236 22600 3288
rect 28600 3236 28652 3288
rect 28674 3236 28726 3288
rect 28748 3236 28800 3288
rect 35893 3238 35945 3290
rect 35957 3238 36009 3290
rect 36021 3238 36073 3290
rect 1353 1846 1469 1962
rect 6202 1846 6318 1962
rect 6350 1846 6466 1962
rect 12102 1846 12218 1962
rect 12250 1846 12366 1962
rect 18002 1846 18118 1962
rect 18150 1846 18266 1962
rect 23902 1846 24018 1962
rect 24050 1846 24166 1962
rect 29802 1846 29918 1962
rect 29950 1846 30066 1962
rect 33230 1846 33346 1962
rect 33374 1846 33490 1962
rect 811 1301 927 1417
rect 34552 1301 34668 1417
rect 7800 -28 7852 24
rect 7874 -28 7926 24
rect 7948 -28 8000 24
rect 14000 -28 14052 24
rect 14074 -28 14126 24
rect 14148 -28 14200 24
rect 22400 -28 22452 24
rect 22474 -28 22526 24
rect 22548 -28 22600 24
rect 28600 -28 28652 24
rect 28674 -28 28726 24
rect 28748 -28 28800 24
rect 35895 -26 35947 26
rect 35959 -26 36011 26
rect 36023 -26 36075 26
<< metal2 >>
rect 7800 7644 8000 7654
rect 7800 7640 7820 7644
rect 7880 7640 7920 7644
rect 7980 7640 8000 7644
rect 7800 7584 7820 7588
rect 7880 7584 7920 7588
rect 7980 7584 8000 7588
rect 7800 7574 8000 7584
rect 3578 6327 3757 6333
rect 2884 6315 3757 6327
rect 2884 6199 3609 6315
rect 3725 6199 3757 6315
rect 2884 6187 3757 6199
rect 2884 4010 3024 6187
rect 3578 6181 3757 6187
rect 9364 5784 9524 7874
rect 14000 7644 14200 7654
rect 14000 7640 14020 7644
rect 14080 7640 14120 7644
rect 14180 7640 14200 7644
rect 14000 7584 14020 7588
rect 14080 7584 14120 7588
rect 14180 7584 14200 7588
rect 14000 7574 14200 7584
rect 15264 5784 15424 7874
rect 21164 5784 21324 7874
rect 22400 7644 22600 7654
rect 22400 7640 22420 7644
rect 22480 7640 22520 7644
rect 22580 7640 22600 7644
rect 22400 7584 22420 7588
rect 22480 7584 22520 7588
rect 22580 7584 22600 7588
rect 22400 7574 22600 7584
rect 27064 5784 27224 7874
rect 28600 7644 28800 7654
rect 28600 7640 28620 7644
rect 28680 7640 28720 7644
rect 28780 7640 28800 7644
rect 28600 7584 28620 7588
rect 28680 7584 28720 7588
rect 28780 7584 28800 7588
rect 28600 7574 28800 7584
rect 34488 7642 34688 7674
rect 34488 7590 34498 7642
rect 34550 7590 34562 7642
rect 34614 7590 34626 7642
rect 34678 7590 34688 7642
rect 32894 6327 33078 6333
rect 32894 6315 33898 6327
rect 32894 6199 32896 6315
rect 33076 6199 33898 6315
rect 32894 6187 33898 6199
rect 32894 6181 33078 6187
rect 800 3870 3024 4010
rect 3424 5770 3773 5782
rect 3424 5654 3585 5770
rect 3765 5654 3773 5770
rect 3424 5642 3773 5654
rect 9310 5770 9578 5784
rect 9310 5654 9312 5770
rect 9428 5654 9460 5770
rect 9576 5654 9578 5770
rect 9310 5642 9578 5654
rect 15210 5770 15478 5784
rect 15210 5654 15212 5770
rect 15328 5654 15360 5770
rect 15476 5654 15478 5770
rect 15210 5642 15478 5654
rect 21110 5770 21378 5784
rect 21110 5654 21112 5770
rect 21228 5654 21260 5770
rect 21376 5654 21378 5770
rect 21110 5642 21378 5654
rect 27010 5770 27278 5784
rect 27010 5654 27012 5770
rect 27128 5654 27160 5770
rect 27276 5654 27278 5770
rect 27010 5642 27278 5654
rect 32890 5770 33358 5782
rect 32890 5654 32894 5770
rect 33074 5654 33358 5770
rect 32890 5642 33358 5654
rect 800 3707 940 3870
rect 799 2593 940 3707
rect 3424 3470 3564 5642
rect 7800 4380 8000 4390
rect 7800 4376 7820 4380
rect 7880 4376 7920 4380
rect 7980 4376 8000 4380
rect 7800 4320 7820 4324
rect 7880 4320 7920 4324
rect 7980 4320 8000 4324
rect 7800 4310 8000 4320
rect 14000 4380 14200 4390
rect 14000 4376 14020 4380
rect 14080 4376 14120 4380
rect 14180 4376 14200 4380
rect 14000 4320 14020 4324
rect 14080 4320 14120 4324
rect 14180 4320 14200 4324
rect 14000 4310 14200 4320
rect 22400 4380 22600 4390
rect 22400 4376 22420 4380
rect 22480 4376 22520 4380
rect 22580 4376 22600 4380
rect 22400 4320 22420 4324
rect 22480 4320 22520 4324
rect 22580 4320 22600 4324
rect 22400 4310 22600 4320
rect 28600 4380 28800 4390
rect 28600 4376 28620 4380
rect 28680 4376 28720 4380
rect 28780 4376 28800 4380
rect 28600 4320 28620 4324
rect 28680 4320 28720 4324
rect 28780 4320 28800 4324
rect 28600 4310 28800 4320
rect 1341 3330 3564 3470
rect 799 1417 939 2593
rect 1341 1962 1481 3330
rect 1341 1846 1353 1962
rect 1469 1846 1481 1962
rect 1341 1834 1481 1846
rect 799 1301 811 1417
rect 927 1301 939 1417
rect 799 1283 939 1301
rect 2654 -258 2814 3330
rect 7800 3292 8000 3302
rect 7800 3288 7820 3292
rect 7880 3288 7920 3292
rect 7980 3288 8000 3292
rect 7800 3232 7820 3236
rect 7880 3232 7920 3236
rect 7980 3232 8000 3236
rect 7800 3222 8000 3232
rect 14000 3292 14200 3302
rect 14000 3288 14020 3292
rect 14080 3288 14120 3292
rect 14180 3288 14200 3292
rect 14000 3232 14020 3236
rect 14080 3232 14120 3236
rect 14180 3232 14200 3236
rect 14000 3222 14200 3232
rect 22400 3292 22600 3302
rect 22400 3288 22420 3292
rect 22480 3288 22520 3292
rect 22580 3288 22600 3292
rect 22400 3232 22420 3236
rect 22480 3232 22520 3236
rect 22580 3232 22600 3236
rect 22400 3222 22600 3232
rect 28600 3292 28800 3302
rect 28600 3288 28620 3292
rect 28680 3288 28720 3292
rect 28780 3288 28800 3292
rect 28600 3232 28620 3236
rect 28680 3232 28720 3236
rect 28780 3232 28800 3236
rect 28600 3222 28800 3232
rect 33218 1974 33358 5642
rect 33758 3527 33898 6187
rect 34488 4448 34688 7590
rect 34488 4382 36700 4448
rect 34488 4330 34631 4382
rect 34683 4330 34706 4382
rect 34758 4330 34782 4382
rect 34834 4330 34857 4382
rect 34909 4330 34932 4382
rect 34984 4330 35007 4382
rect 35059 4330 35083 4382
rect 35135 4330 35158 4382
rect 35210 4330 35233 4382
rect 35285 4330 35307 4382
rect 35359 4330 35383 4382
rect 35435 4330 36700 4382
rect 34488 4288 36700 4330
rect 34488 4248 36088 4288
rect 35888 4140 36087 4248
rect 35888 3900 36088 4140
rect 35888 3820 35950 3900
rect 36030 3820 36088 3900
rect 35888 3794 36088 3820
rect 35888 3714 35950 3794
rect 36030 3714 36088 3794
rect 33758 3387 34680 3527
rect 6200 1962 6468 1974
rect 6200 1846 6202 1962
rect 6318 1846 6350 1962
rect 6466 1846 6468 1962
rect 6200 1838 6468 1846
rect 12100 1962 12368 1974
rect 12100 1846 12102 1962
rect 12218 1846 12250 1962
rect 12366 1846 12368 1962
rect 12100 1838 12368 1846
rect 18000 1962 18268 1974
rect 18000 1846 18002 1962
rect 18118 1846 18150 1962
rect 18266 1846 18268 1962
rect 18000 1838 18268 1846
rect 23900 1962 24168 1974
rect 23900 1846 23902 1962
rect 24018 1846 24050 1962
rect 24166 1846 24168 1962
rect 23900 1838 24168 1846
rect 29800 1962 30068 1974
rect 29800 1846 29802 1962
rect 29918 1846 29950 1962
rect 30066 1846 30068 1962
rect 29800 1838 30068 1846
rect 33218 1962 33492 1974
rect 33218 1846 33230 1962
rect 33346 1846 33374 1962
rect 33490 1846 33492 1962
rect 6254 -258 6414 1838
rect 7800 28 8000 38
rect 7800 24 7820 28
rect 7880 24 7920 28
rect 7980 24 8000 28
rect 7800 -32 7820 -28
rect 7880 -32 7920 -28
rect 7980 -32 8000 -28
rect 7800 -42 8000 -32
rect 12154 -258 12314 1838
rect 14000 28 14200 38
rect 14000 24 14020 28
rect 14080 24 14120 28
rect 14180 24 14200 28
rect 14000 -32 14020 -28
rect 14080 -32 14120 -28
rect 14180 -32 14200 -28
rect 14000 -42 14200 -32
rect 18054 -258 18214 1838
rect 22400 28 22600 38
rect 22400 24 22420 28
rect 22480 24 22520 28
rect 22580 24 22600 28
rect 22400 -32 22420 -28
rect 22480 -32 22520 -28
rect 22580 -32 22600 -28
rect 22400 -42 22600 -32
rect 23954 -258 24114 1838
rect 28600 28 28800 38
rect 28600 24 28620 28
rect 28680 24 28720 28
rect 28780 24 28800 28
rect 28600 -32 28620 -28
rect 28680 -32 28720 -28
rect 28780 -32 28800 -28
rect 28600 -42 28800 -32
rect 29854 -258 30014 1838
rect 33218 1828 33492 1846
rect 33272 -258 33432 1828
rect 34540 1417 34680 3387
rect 34540 1301 34552 1417
rect 34668 1301 34680 1417
rect 34540 1289 34680 1301
rect 35888 3290 36088 3714
rect 35888 3238 35893 3290
rect 35945 3238 35957 3290
rect 36009 3238 36021 3290
rect 36073 3238 36088 3290
rect 35888 26 36088 3238
rect 35888 -26 35895 26
rect 35947 -26 35959 26
rect 36011 -26 36023 26
rect 36075 -26 36088 26
rect 35888 -58 36088 -26
<< via2 >>
rect 7820 7640 7880 7644
rect 7920 7640 7980 7644
rect 7820 7588 7852 7640
rect 7852 7588 7874 7640
rect 7874 7588 7880 7640
rect 7920 7588 7926 7640
rect 7926 7588 7948 7640
rect 7948 7588 7980 7640
rect 7820 7584 7880 7588
rect 7920 7584 7980 7588
rect 14020 7640 14080 7644
rect 14120 7640 14180 7644
rect 14020 7588 14052 7640
rect 14052 7588 14074 7640
rect 14074 7588 14080 7640
rect 14120 7588 14126 7640
rect 14126 7588 14148 7640
rect 14148 7588 14180 7640
rect 14020 7584 14080 7588
rect 14120 7584 14180 7588
rect 22420 7640 22480 7644
rect 22520 7640 22580 7644
rect 22420 7588 22452 7640
rect 22452 7588 22474 7640
rect 22474 7588 22480 7640
rect 22520 7588 22526 7640
rect 22526 7588 22548 7640
rect 22548 7588 22580 7640
rect 22420 7584 22480 7588
rect 22520 7584 22580 7588
rect 28620 7640 28680 7644
rect 28720 7640 28780 7644
rect 28620 7588 28652 7640
rect 28652 7588 28674 7640
rect 28674 7588 28680 7640
rect 28720 7588 28726 7640
rect 28726 7588 28748 7640
rect 28748 7588 28780 7640
rect 28620 7584 28680 7588
rect 28720 7584 28780 7588
rect 7820 4376 7880 4380
rect 7920 4376 7980 4380
rect 7820 4324 7852 4376
rect 7852 4324 7874 4376
rect 7874 4324 7880 4376
rect 7920 4324 7926 4376
rect 7926 4324 7948 4376
rect 7948 4324 7980 4376
rect 7820 4320 7880 4324
rect 7920 4320 7980 4324
rect 14020 4376 14080 4380
rect 14120 4376 14180 4380
rect 14020 4324 14052 4376
rect 14052 4324 14074 4376
rect 14074 4324 14080 4376
rect 14120 4324 14126 4376
rect 14126 4324 14148 4376
rect 14148 4324 14180 4376
rect 14020 4320 14080 4324
rect 14120 4320 14180 4324
rect 22420 4376 22480 4380
rect 22520 4376 22580 4380
rect 22420 4324 22452 4376
rect 22452 4324 22474 4376
rect 22474 4324 22480 4376
rect 22520 4324 22526 4376
rect 22526 4324 22548 4376
rect 22548 4324 22580 4376
rect 22420 4320 22480 4324
rect 22520 4320 22580 4324
rect 28620 4376 28680 4380
rect 28720 4376 28780 4380
rect 28620 4324 28652 4376
rect 28652 4324 28674 4376
rect 28674 4324 28680 4376
rect 28720 4324 28726 4376
rect 28726 4324 28748 4376
rect 28748 4324 28780 4376
rect 28620 4320 28680 4324
rect 28720 4320 28780 4324
rect 7820 3288 7880 3292
rect 7920 3288 7980 3292
rect 7820 3236 7852 3288
rect 7852 3236 7874 3288
rect 7874 3236 7880 3288
rect 7920 3236 7926 3288
rect 7926 3236 7948 3288
rect 7948 3236 7980 3288
rect 7820 3232 7880 3236
rect 7920 3232 7980 3236
rect 14020 3288 14080 3292
rect 14120 3288 14180 3292
rect 14020 3236 14052 3288
rect 14052 3236 14074 3288
rect 14074 3236 14080 3288
rect 14120 3236 14126 3288
rect 14126 3236 14148 3288
rect 14148 3236 14180 3288
rect 14020 3232 14080 3236
rect 14120 3232 14180 3236
rect 22420 3288 22480 3292
rect 22520 3288 22580 3292
rect 22420 3236 22452 3288
rect 22452 3236 22474 3288
rect 22474 3236 22480 3288
rect 22520 3236 22526 3288
rect 22526 3236 22548 3288
rect 22548 3236 22580 3288
rect 22420 3232 22480 3236
rect 22520 3232 22580 3236
rect 28620 3288 28680 3292
rect 28720 3288 28780 3292
rect 28620 3236 28652 3288
rect 28652 3236 28674 3288
rect 28674 3236 28680 3288
rect 28720 3236 28726 3288
rect 28726 3236 28748 3288
rect 28748 3236 28780 3288
rect 28620 3232 28680 3236
rect 28720 3232 28780 3236
rect 35950 3820 36030 3900
rect 35950 3714 36030 3794
rect 7820 24 7880 28
rect 7920 24 7980 28
rect 7820 -28 7852 24
rect 7852 -28 7874 24
rect 7874 -28 7880 24
rect 7920 -28 7926 24
rect 7926 -28 7948 24
rect 7948 -28 7980 24
rect 7820 -32 7880 -28
rect 7920 -32 7980 -28
rect 14020 24 14080 28
rect 14120 24 14180 28
rect 14020 -28 14052 24
rect 14052 -28 14074 24
rect 14074 -28 14080 24
rect 14120 -28 14126 24
rect 14126 -28 14148 24
rect 14148 -28 14180 24
rect 14020 -32 14080 -28
rect 14120 -32 14180 -28
rect 22420 24 22480 28
rect 22520 24 22580 28
rect 22420 -28 22452 24
rect 22452 -28 22474 24
rect 22474 -28 22480 24
rect 22520 -28 22526 24
rect 22526 -28 22548 24
rect 22548 -28 22580 24
rect 22420 -32 22480 -28
rect 22520 -32 22580 -28
rect 28620 24 28680 28
rect 28720 24 28780 28
rect 28620 -28 28652 24
rect 28652 -28 28674 24
rect 28674 -28 28680 24
rect 28720 -28 28726 24
rect 28726 -28 28748 24
rect 28748 -28 28780 24
rect 28620 -32 28680 -28
rect 28720 -32 28780 -28
<< metal3 >>
rect 7800 7644 8000 7664
rect 7800 7584 7820 7644
rect 7880 7584 7920 7644
rect 7980 7584 8000 7644
rect 7800 4380 8000 7584
rect 7800 4320 7820 4380
rect 7880 4320 7920 4380
rect 7980 4320 8000 4380
rect 7800 3922 8000 4320
rect 14000 7644 14200 7664
rect 14000 7584 14020 7644
rect 14080 7584 14120 7644
rect 14180 7584 14200 7644
rect 14000 4380 14200 7584
rect 14000 4320 14020 4380
rect 14080 4320 14120 4380
rect 14180 4320 14200 4380
rect 14000 3922 14200 4320
rect 22400 7644 22600 7664
rect 22400 7584 22420 7644
rect 22480 7584 22520 7644
rect 22580 7584 22600 7644
rect 22400 4380 22600 7584
rect 22400 4320 22420 4380
rect 22480 4320 22520 4380
rect 22580 4320 22600 4380
rect 22400 3922 22600 4320
rect 28600 7644 28800 7664
rect 28600 7584 28620 7644
rect 28680 7584 28720 7644
rect 28780 7584 28800 7644
rect 28600 4380 28800 7584
rect 28600 4320 28620 4380
rect 28680 4320 28720 4380
rect 28780 4320 28800 4380
rect 28600 3922 28800 4320
rect 7800 3900 36088 3922
rect 7800 3820 35950 3900
rect 36030 3820 36088 3900
rect 7800 3794 36088 3820
rect 7800 3714 35950 3794
rect 36030 3714 36088 3794
rect 7800 3692 36088 3714
rect 7800 3292 8000 3692
rect 7800 3232 7820 3292
rect 7880 3232 7920 3292
rect 7980 3232 8000 3292
rect 7800 28 8000 3232
rect 7800 -32 7820 28
rect 7880 -32 7920 28
rect 7980 -32 8000 28
rect 7800 -48 8000 -32
rect 14000 3292 14200 3692
rect 14000 3232 14020 3292
rect 14080 3232 14120 3292
rect 14180 3232 14200 3292
rect 14000 28 14200 3232
rect 14000 -32 14020 28
rect 14080 -32 14120 28
rect 14180 -32 14200 28
rect 14000 -48 14200 -32
rect 22400 3292 22600 3692
rect 22400 3232 22420 3292
rect 22480 3232 22520 3292
rect 22580 3232 22600 3292
rect 22400 28 22600 3232
rect 22400 -32 22420 28
rect 22480 -32 22520 28
rect 22580 -32 22600 28
rect 22400 -48 22600 -32
rect 28600 3292 28800 3692
rect 28600 3232 28620 3292
rect 28680 3232 28720 3292
rect 28780 3232 28800 3292
rect 28600 28 28800 3232
rect 28600 -32 28620 28
rect 28680 -32 28720 28
rect 28780 -32 28800 28
rect 28600 -48 28800 -32
use inv_ver_3-1  inv_ver_3-1_0
timestamp 1622803027
transform -1 0 6300 0 1 -48
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_1
timestamp 1622803027
transform -1 0 12200 0 1 -48
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_2
timestamp 1622803027
transform -1 0 18100 0 1 -48
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_3
timestamp 1622803027
transform -1 0 24000 0 1 -48
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_4
timestamp 1622803027
transform -1 0 29900 0 1 -48
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_5
timestamp 1622803027
transform -1 0 35800 0 1 -48
box 0 -10 5900 3372
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag/
timestamp 1621367673
transform 1 0 764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag/
timestamp 1621367673
transform 1 0 1598 0 1 5440
box -38 -48 314 592
use inv_ver_3-1  inv_ver_3-1_6
timestamp 1622803027
transform 1 0 3578 0 -1 7664
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_7
timestamp 1622803027
transform 1 0 9478 0 -1 7664
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_8
timestamp 1622803027
transform 1 0 15378 0 -1 7664
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_9
timestamp 1622803027
transform 1 0 21278 0 -1 7664
box 0 -10 5900 3372
use inv_ver_3-1  inv_ver_3-1_10
timestamp 1622803027
transform 1 0 27178 0 -1 7664
box 0 -10 5900 3372
<< labels >>
flabel metal1 s 0 5392 400 5488 1 FreeSans 2343 0 0 0 vssd1
flabel metal1 s 3200 7024 3600 7120 1 FreeSans 2343 0 0 0 vccd1
flabel metal1 s 3001 4848 3401 4944 1 FreeSans 2343 0 0 0 vccd1
flabel metal1 s 3658 5936 4058 6032 5 FreeSans 2343 180 0 0 vccd1
flabel metal2 s 27064 7674 27224 7874 1 FreeSans 2343 0 0 0 p[9]
flabel metal2 s 21164 7674 21324 7874 1 FreeSans 2343 0 0 0 p[8]
flabel metal2 s 15264 7674 15424 7874 1 FreeSans 2343 0 0 0 p[7]
flabel metal2 s 9364 7674 9524 7874 1 FreeSans 2343 0 0 0 p[6]
flabel metal1 s 27044 6192 27342 6320 1 FreeSans 2343 0 0 0 pn_9
flabel metal1 s 21152 6192 21450 6320 1 FreeSans 2343 0 0 0 pn_8
flabel metal1 s 15248 6194 15546 6322 1 FreeSans 2343 0 0 0 pn_7
flabel metal1 s 9336 6192 9634 6320 1 FreeSans 2343 0 0 0 pn_6
flabel metal2 s 33272 -258 33432 -58 1 FreeSans 2343 0 0 0 p[10]
flabel metal2 s 2654 -258 2814 -58 1 FreeSans 2343 0 0 0 p[5]
flabel metal2 s 6254 -258 6414 -58 1 FreeSans 2343 0 0 0 p[4]
flabel metal2 s 12154 -258 12314 -58 1 FreeSans 2343 0 0 0 p[3]
flabel metal2 s 18054 -258 18214 -58 1 FreeSans 2343 0 0 0 p[2]
flabel metal2 s 23954 -258 24114 -58 1 FreeSans 2343 0 0 0 p[1]
flabel metal2 s 29854 -258 30014 -58 1 FreeSans 2343 0 0 0 p[0]
flabel metal1 s 0 2672 400 2768 1 FreeSans 2343 0 0 0 vccd1
flabel metal1 s 0 496 400 592 1 FreeSans 2343 0 0 0 vccd1
flabel metal2 s 34364 3388 34680 3526 1 FreeSans 2343 0 0 0 pn_10
flabel metal2 s 800 3872 1116 4010 1 FreeSans 2343 0 0 0 pn_5
flabel metal1 s 6144 1296 6442 1424 1 FreeSans 2343 180 0 0 pn_4
flabel metal1 s 12044 1294 12342 1422 1 FreeSans 2343 0 0 0 pn_3
flabel metal1 s 17956 1294 18254 1422 1 FreeSans 2343 0 0 0 pn_2
flabel metal1 s 23852 1294 24150 1422 1 FreeSans 2343 0 0 0 pn_1
flabel metal1 s 29768 1294 30052 1424 1 FreeSans 2343 0 0 0 pn_0
flabel locali 1326 5815 1496 5875 1 FreeSans 400 0 0 0 hi_logic
flabel locali 807 5652 857 5685 1 FreeSans 400 0 0 0 enb
flabel metal3 32038 3692 32700 3922 1 FreeSans 2 0 0 0 v_crt
flabel metal2 s 36500 4288 36700 4448 1 FreeSans 2343 0 0 0 input_analog
<< end >>
